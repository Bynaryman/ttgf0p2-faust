module process(
  input [7:0] in0,
  input  in0_valid,
  input  start_valid,
  input  clk,
  input  rst,
  input  out0_ready,
  input  end_ready,
  output  in0_ready,
  output  start_ready,
  output [7:0] out0,
  output  out0_valid,
  output  end_valid
);
  wire  fork0_outs_0_valid;
  wire  fork0_outs_0_ready;
  wire  fork0_outs_1_valid;
  wire  fork0_outs_1_ready;
  wire  fork0_outs_2_valid;
  wire  fork0_outs_2_ready;
  wire  fork0_outs_3_valid;
  wire  fork0_outs_3_ready;
  wire  fork0_outs_4_valid;
  wire  fork0_outs_4_ready;
  wire  fork0_outs_5_valid;
  wire  fork0_outs_5_ready;
  wire  fork0_outs_6_valid;
  wire  fork0_outs_6_ready;
  wire  fork0_outs_7_valid;
  wire  fork0_outs_7_ready;
  wire  fork0_outs_8_valid;
  wire  fork0_outs_8_ready;
  wire  fork0_outs_9_valid;
  wire  fork0_outs_9_ready;
  wire  fork0_outs_10_valid;
  wire  fork0_outs_10_ready;
  wire  fork0_outs_11_valid;
  wire  fork0_outs_11_ready;
  wire  fork0_outs_12_valid;
  wire  fork0_outs_12_ready;
  wire [7:0] fork1_outs_0;
  wire  fork1_outs_0_valid;
  wire  fork1_outs_0_ready;
  wire [7:0] fork1_outs_1;
  wire  fork1_outs_1_valid;
  wire  fork1_outs_1_ready;
  wire [4:0] trunci23_outs;
  wire  trunci23_outs_valid;
  wire  trunci23_outs_ready;
  wire  source0_outs_valid;
  wire  source0_outs_ready;
  wire [0:0] constant212_outs;
  wire  constant212_outs_valid;
  wire  constant212_outs_ready;
  wire [2:0] extsi99_outs;
  wire  extsi99_outs_valid;
  wire  extsi99_outs_ready;
  wire [7:0] constant94_outs;
  wire  constant94_outs_valid;
  wire  constant94_outs_ready;
  wire [6:0] constant213_outs;
  wire  constant213_outs_valid;
  wire  constant213_outs_ready;
  wire [11:0] constant96_outs;
  wire  constant96_outs_valid;
  wire  constant96_outs_ready;
  wire [13:0] constant97_outs;
  wire  constant97_outs_valid;
  wire  constant97_outs_ready;
  wire [17:0] constant98_outs;
  wire  constant98_outs_valid;
  wire  constant98_outs_ready;
  wire [20:0] constant99_outs;
  wire  constant99_outs_valid;
  wire  constant99_outs_ready;
  wire [23:0] constant100_outs;
  wire  constant100_outs_valid;
  wire  constant100_outs_ready;
  wire [26:0] constant101_outs;
  wire  constant101_outs_valid;
  wire  constant101_outs_ready;
  wire [29:0] constant102_outs;
  wire  constant102_outs_valid;
  wire  constant102_outs_ready;
  wire [33:0] constant103_outs;
  wire  constant103_outs_valid;
  wire  constant103_outs_ready;
  wire [33:0] constant214_outs;
  wire  constant214_outs_valid;
  wire  constant214_outs_ready;
  wire  source1_outs_valid;
  wire  source1_outs_ready;
  wire [3:0] constant215_outs;
  wire  constant215_outs_valid;
  wire  constant215_outs_ready;
  wire [7:0] extsi43_outs;
  wire  extsi43_outs_valid;
  wire  extsi43_outs_ready;
  wire [7:0] shrui0_result;
  wire  shrui0_result_valid;
  wire  shrui0_result_ready;
  wire [2:0] trunci0_outs;
  wire  trunci0_outs_valid;
  wire  trunci0_outs_ready;
  wire [2:0] fork2_outs_0;
  wire  fork2_outs_0_valid;
  wire  fork2_outs_0_ready;
  wire [2:0] fork2_outs_1;
  wire  fork2_outs_1_valid;
  wire  fork2_outs_1_ready;
  wire [0:0] cmpi0_result;
  wire  cmpi0_result_valid;
  wire  cmpi0_result_ready;
  wire [0:0] fork3_outs_0;
  wire  fork3_outs_0_valid;
  wire  fork3_outs_0_ready;
  wire [0:0] fork3_outs_1;
  wire  fork3_outs_1_valid;
  wire  fork3_outs_1_ready;
  wire [0:0] fork3_outs_2;
  wire  fork3_outs_2_valid;
  wire  fork3_outs_2_ready;
  wire [0:0] fork3_outs_3;
  wire  fork3_outs_3_valid;
  wire  fork3_outs_3_ready;
  wire [0:0] fork3_outs_4;
  wire  fork3_outs_4_valid;
  wire  fork3_outs_4_ready;
  wire [0:0] fork3_outs_5;
  wire  fork3_outs_5_valid;
  wire  fork3_outs_5_ready;
  wire [0:0] fork3_outs_6;
  wire  fork3_outs_6_valid;
  wire  fork3_outs_6_ready;
  wire [0:0] fork3_outs_7;
  wire  fork3_outs_7_valid;
  wire  fork3_outs_7_ready;
  wire [0:0] fork3_outs_8;
  wire  fork3_outs_8_valid;
  wire  fork3_outs_8_ready;
  wire [0:0] fork3_outs_9;
  wire  fork3_outs_9_valid;
  wire  fork3_outs_9_ready;
  wire [0:0] fork3_outs_10;
  wire  fork3_outs_10_valid;
  wire  fork3_outs_10_ready;
  wire [0:0] fork3_outs_11;
  wire  fork3_outs_11_valid;
  wire  fork3_outs_11_ready;
  wire [0:0] fork3_outs_12;
  wire  fork3_outs_12_valid;
  wire  fork3_outs_12_ready;
  wire [0:0] fork3_outs_13;
  wire  fork3_outs_13_valid;
  wire  fork3_outs_13_ready;
  wire [33:0] cond_br8_trueOut;
  wire  cond_br8_trueOut_valid;
  wire  cond_br8_trueOut_ready;
  wire [33:0] cond_br8_falseOut;
  wire  cond_br8_falseOut_valid;
  wire  cond_br8_falseOut_ready;
  wire [35:0] extsi100_outs;
  wire  extsi100_outs_valid;
  wire  extsi100_outs_ready;
  wire [33:0] cond_br9_trueOut;
  wire  cond_br9_trueOut_valid;
  wire  cond_br9_trueOut_ready;
  wire [33:0] cond_br9_falseOut;
  wire  cond_br9_falseOut_valid;
  wire  cond_br9_falseOut_ready;
  wire [29:0] cond_br10_trueOut;
  wire  cond_br10_trueOut_valid;
  wire  cond_br10_trueOut_ready;
  wire [29:0] cond_br10_falseOut;
  wire  cond_br10_falseOut_valid;
  wire  cond_br10_falseOut_ready;
  wire [26:0] cond_br11_trueOut;
  wire  cond_br11_trueOut_valid;
  wire  cond_br11_trueOut_ready;
  wire [26:0] cond_br11_falseOut;
  wire  cond_br11_falseOut_valid;
  wire  cond_br11_falseOut_ready;
  wire [23:0] cond_br12_trueOut;
  wire  cond_br12_trueOut_valid;
  wire  cond_br12_trueOut_ready;
  wire [23:0] cond_br12_falseOut;
  wire  cond_br12_falseOut_valid;
  wire  cond_br12_falseOut_ready;
  wire [20:0] cond_br13_trueOut;
  wire  cond_br13_trueOut_valid;
  wire  cond_br13_trueOut_ready;
  wire [20:0] cond_br13_falseOut;
  wire  cond_br13_falseOut_valid;
  wire  cond_br13_falseOut_ready;
  wire [17:0] cond_br14_trueOut;
  wire  cond_br14_trueOut_valid;
  wire  cond_br14_trueOut_ready;
  wire [17:0] cond_br14_falseOut;
  wire  cond_br14_falseOut_valid;
  wire  cond_br14_falseOut_ready;
  wire [13:0] cond_br15_trueOut;
  wire  cond_br15_trueOut_valid;
  wire  cond_br15_trueOut_ready;
  wire [13:0] cond_br15_falseOut;
  wire  cond_br15_falseOut_valid;
  wire  cond_br15_falseOut_ready;
  wire [11:0] cond_br16_trueOut;
  wire  cond_br16_trueOut_valid;
  wire  cond_br16_trueOut_ready;
  wire [11:0] cond_br16_falseOut;
  wire  cond_br16_falseOut_valid;
  wire  cond_br16_falseOut_ready;
  wire [6:0] cond_br17_trueOut;
  wire  cond_br17_trueOut_valid;
  wire  cond_br17_trueOut_ready;
  wire [6:0] cond_br17_falseOut;
  wire  cond_br17_falseOut_valid;
  wire  cond_br17_falseOut_ready;
  wire [7:0] extsi101_outs;
  wire  extsi101_outs_valid;
  wire  extsi101_outs_ready;
  wire [7:0] cond_br18_trueOut;
  wire  cond_br18_trueOut_valid;
  wire  cond_br18_trueOut_ready;
  wire [7:0] cond_br18_falseOut;
  wire  cond_br18_falseOut_valid;
  wire  cond_br18_falseOut_ready;
  wire [4:0] cond_br19_trueOut;
  wire  cond_br19_trueOut_valid;
  wire  cond_br19_trueOut_ready;
  wire [4:0] cond_br19_falseOut;
  wire  cond_br19_falseOut_valid;
  wire  cond_br19_falseOut_ready;
  wire  cond_br20_trueOut_valid;
  wire  cond_br20_trueOut_ready;
  wire  cond_br20_falseOut_valid;
  wire  cond_br20_falseOut_ready;
  wire [2:0] cond_br21_trueOut;
  wire  cond_br21_trueOut_valid;
  wire  cond_br21_trueOut_ready;
  wire [2:0] cond_br21_falseOut;
  wire  cond_br21_falseOut_valid;
  wire  cond_br21_falseOut_ready;
  wire [2:0] buffer2_outs;
  wire  buffer2_outs_valid;
  wire  buffer2_outs_ready;
  wire [2:0] buffer3_outs;
  wire  buffer3_outs_valid;
  wire  buffer3_outs_ready;
  wire [2:0] fork4_outs_0;
  wire  fork4_outs_0_valid;
  wire  fork4_outs_0_ready;
  wire [2:0] fork4_outs_1;
  wire  fork4_outs_1_valid;
  wire  fork4_outs_1_ready;
  wire  buffer4_outs_valid;
  wire  buffer4_outs_ready;
  wire  buffer5_outs_valid;
  wire  buffer5_outs_ready;
  wire  fork5_outs_0_valid;
  wire  fork5_outs_0_ready;
  wire  fork5_outs_1_valid;
  wire  fork5_outs_1_ready;
  wire  fork5_outs_2_valid;
  wire  fork5_outs_2_ready;
  wire  fork5_outs_3_valid;
  wire  fork5_outs_3_ready;
  wire  fork5_outs_4_valid;
  wire  fork5_outs_4_ready;
  wire  fork5_outs_5_valid;
  wire  fork5_outs_5_ready;
  wire  fork5_outs_6_valid;
  wire  fork5_outs_6_ready;
  wire  fork5_outs_7_valid;
  wire  fork5_outs_7_ready;
  wire  fork5_outs_8_valid;
  wire  fork5_outs_8_ready;
  wire  fork5_outs_9_valid;
  wire  fork5_outs_9_ready;
  wire  fork5_outs_10_valid;
  wire  fork5_outs_10_ready;
  wire  fork5_outs_11_valid;
  wire  fork5_outs_11_ready;
  wire [34:0] constant216_outs;
  wire  constant216_outs_valid;
  wire  constant216_outs_ready;
  wire [32:0] constant217_outs;
  wire  constant217_outs_valid;
  wire  constant217_outs_ready;
  wire [29:0] constant108_outs;
  wire  constant108_outs_valid;
  wire  constant108_outs_ready;
  wire [26:0] constant109_outs;
  wire  constant109_outs_valid;
  wire  constant109_outs_ready;
  wire [23:0] constant110_outs;
  wire  constant110_outs_valid;
  wire  constant110_outs_ready;
  wire [20:0] constant111_outs;
  wire  constant111_outs_valid;
  wire  constant111_outs_ready;
  wire [17:0] constant112_outs;
  wire  constant112_outs_valid;
  wire  constant112_outs_ready;
  wire [13:0] constant113_outs;
  wire  constant113_outs_valid;
  wire  constant113_outs_ready;
  wire [8:0] constant218_outs;
  wire  constant218_outs_valid;
  wire  constant218_outs_ready;
  wire [7:0] constant115_outs;
  wire  constant115_outs_valid;
  wire  constant115_outs_ready;
  wire [7:0] constant116_outs;
  wire  constant116_outs_valid;
  wire  constant116_outs_ready;
  wire  source2_outs_valid;
  wire  source2_outs_ready;
  wire [1:0] constant219_outs;
  wire  constant219_outs_valid;
  wire  constant219_outs_ready;
  wire [2:0] extsi102_outs;
  wire  extsi102_outs_valid;
  wire  extsi102_outs_ready;
  wire [0:0] cmpi1_result;
  wire  cmpi1_result_valid;
  wire  cmpi1_result_ready;
  wire [0:0] fork6_outs_0;
  wire  fork6_outs_0_valid;
  wire  fork6_outs_0_ready;
  wire [0:0] fork6_outs_1;
  wire  fork6_outs_1_valid;
  wire  fork6_outs_1_ready;
  wire [0:0] fork6_outs_2;
  wire  fork6_outs_2_valid;
  wire  fork6_outs_2_ready;
  wire [0:0] fork6_outs_3;
  wire  fork6_outs_3_valid;
  wire  fork6_outs_3_ready;
  wire [0:0] fork6_outs_4;
  wire  fork6_outs_4_valid;
  wire  fork6_outs_4_ready;
  wire [0:0] fork6_outs_5;
  wire  fork6_outs_5_valid;
  wire  fork6_outs_5_ready;
  wire [0:0] fork6_outs_6;
  wire  fork6_outs_6_valid;
  wire  fork6_outs_6_ready;
  wire [0:0] fork6_outs_7;
  wire  fork6_outs_7_valid;
  wire  fork6_outs_7_ready;
  wire [0:0] fork6_outs_8;
  wire  fork6_outs_8_valid;
  wire  fork6_outs_8_ready;
  wire [0:0] fork6_outs_9;
  wire  fork6_outs_9_valid;
  wire  fork6_outs_9_ready;
  wire [0:0] fork6_outs_10;
  wire  fork6_outs_10_valid;
  wire  fork6_outs_10_ready;
  wire [0:0] fork6_outs_11;
  wire  fork6_outs_11_valid;
  wire  fork6_outs_11_ready;
  wire [0:0] fork6_outs_12;
  wire  fork6_outs_12_valid;
  wire  fork6_outs_12_ready;
  wire [0:0] fork6_outs_13;
  wire  fork6_outs_13_valid;
  wire  fork6_outs_13_ready;
  wire [34:0] cond_br22_trueOut;
  wire  cond_br22_trueOut_valid;
  wire  cond_br22_trueOut_ready;
  wire [34:0] cond_br22_falseOut;
  wire  cond_br22_falseOut_valid;
  wire  cond_br22_falseOut_ready;
  wire [35:0] extsi103_outs;
  wire  extsi103_outs_valid;
  wire  extsi103_outs_ready;
  wire [32:0] cond_br23_trueOut;
  wire  cond_br23_trueOut_valid;
  wire  cond_br23_trueOut_ready;
  wire [32:0] cond_br23_falseOut;
  wire  cond_br23_falseOut_valid;
  wire  cond_br23_falseOut_ready;
  wire [33:0] extsi104_outs;
  wire  extsi104_outs_valid;
  wire  extsi104_outs_ready;
  wire [29:0] cond_br24_trueOut;
  wire  cond_br24_trueOut_valid;
  wire  cond_br24_trueOut_ready;
  wire [29:0] cond_br24_falseOut;
  wire  cond_br24_falseOut_valid;
  wire  cond_br24_falseOut_ready;
  wire [26:0] cond_br25_trueOut;
  wire  cond_br25_trueOut_valid;
  wire  cond_br25_trueOut_ready;
  wire [26:0] cond_br25_falseOut;
  wire  cond_br25_falseOut_valid;
  wire  cond_br25_falseOut_ready;
  wire [23:0] cond_br26_trueOut;
  wire  cond_br26_trueOut_valid;
  wire  cond_br26_trueOut_ready;
  wire [23:0] cond_br26_falseOut;
  wire  cond_br26_falseOut_valid;
  wire  cond_br26_falseOut_ready;
  wire [20:0] cond_br27_trueOut;
  wire  cond_br27_trueOut_valid;
  wire  cond_br27_trueOut_ready;
  wire [20:0] cond_br27_falseOut;
  wire  cond_br27_falseOut_valid;
  wire  cond_br27_falseOut_ready;
  wire [17:0] cond_br28_trueOut;
  wire  cond_br28_trueOut_valid;
  wire  cond_br28_trueOut_ready;
  wire [17:0] cond_br28_falseOut;
  wire  cond_br28_falseOut_valid;
  wire  cond_br28_falseOut_ready;
  wire [13:0] cond_br29_trueOut;
  wire  cond_br29_trueOut_valid;
  wire  cond_br29_trueOut_ready;
  wire [13:0] cond_br29_falseOut;
  wire  cond_br29_falseOut_valid;
  wire  cond_br29_falseOut_ready;
  wire [8:0] cond_br30_trueOut;
  wire  cond_br30_trueOut_valid;
  wire  cond_br30_trueOut_ready;
  wire [8:0] cond_br30_falseOut;
  wire  cond_br30_falseOut_valid;
  wire  cond_br30_falseOut_ready;
  wire [11:0] extsi105_outs;
  wire  extsi105_outs_valid;
  wire  extsi105_outs_ready;
  wire [7:0] cond_br31_trueOut;
  wire  cond_br31_trueOut_valid;
  wire  cond_br31_trueOut_ready;
  wire [7:0] cond_br31_falseOut;
  wire  cond_br31_falseOut_valid;
  wire  cond_br31_falseOut_ready;
  wire [7:0] cond_br32_trueOut;
  wire  cond_br32_trueOut_valid;
  wire  cond_br32_trueOut_ready;
  wire [7:0] cond_br32_falseOut;
  wire  cond_br32_falseOut_valid;
  wire  cond_br32_falseOut_ready;
  wire [4:0] buffer0_outs;
  wire  buffer0_outs_valid;
  wire  buffer0_outs_ready;
  wire [4:0] buffer1_outs;
  wire  buffer1_outs_valid;
  wire  buffer1_outs_ready;
  wire [4:0] cond_br33_trueOut;
  wire  cond_br33_trueOut_valid;
  wire  cond_br33_trueOut_ready;
  wire [4:0] cond_br33_falseOut;
  wire  cond_br33_falseOut_valid;
  wire  cond_br33_falseOut_ready;
  wire  cond_br34_trueOut_valid;
  wire  cond_br34_trueOut_ready;
  wire  cond_br34_falseOut_valid;
  wire  cond_br34_falseOut_ready;
  wire [2:0] cond_br35_trueOut;
  wire  cond_br35_trueOut_valid;
  wire  cond_br35_trueOut_ready;
  wire [2:0] cond_br35_falseOut;
  wire  cond_br35_falseOut_valid;
  wire  cond_br35_falseOut_ready;
  wire [2:0] buffer8_outs;
  wire  buffer8_outs_valid;
  wire  buffer8_outs_ready;
  wire [2:0] buffer9_outs;
  wire  buffer9_outs_valid;
  wire  buffer9_outs_ready;
  wire [2:0] fork7_outs_0;
  wire  fork7_outs_0_valid;
  wire  fork7_outs_0_ready;
  wire [2:0] fork7_outs_1;
  wire  fork7_outs_1_valid;
  wire  fork7_outs_1_ready;
  wire  buffer10_outs_valid;
  wire  buffer10_outs_ready;
  wire  buffer11_outs_valid;
  wire  buffer11_outs_ready;
  wire  fork8_outs_0_valid;
  wire  fork8_outs_0_ready;
  wire  fork8_outs_1_valid;
  wire  fork8_outs_1_ready;
  wire  fork8_outs_2_valid;
  wire  fork8_outs_2_ready;
  wire  fork8_outs_3_valid;
  wire  fork8_outs_3_ready;
  wire  fork8_outs_4_valid;
  wire  fork8_outs_4_ready;
  wire  fork8_outs_5_valid;
  wire  fork8_outs_5_ready;
  wire  fork8_outs_6_valid;
  wire  fork8_outs_6_ready;
  wire  fork8_outs_7_valid;
  wire  fork8_outs_7_ready;
  wire  fork8_outs_8_valid;
  wire  fork8_outs_8_ready;
  wire  fork8_outs_9_valid;
  wire  fork8_outs_9_ready;
  wire  fork8_outs_10_valid;
  wire  fork8_outs_10_ready;
  wire  fork8_outs_11_valid;
  wire  fork8_outs_11_ready;
  wire [35:0] constant118_outs;
  wire  constant118_outs_valid;
  wire  constant118_outs_ready;
  wire [32:0] constant220_outs;
  wire  constant220_outs_valid;
  wire  constant220_outs_ready;
  wire [29:0] constant120_outs;
  wire  constant120_outs_valid;
  wire  constant120_outs_ready;
  wire [25:0] constant221_outs;
  wire  constant221_outs_valid;
  wire  constant221_outs_ready;
  wire [21:0] constant222_outs;
  wire  constant222_outs_valid;
  wire  constant222_outs_ready;
  wire [20:0] constant123_outs;
  wire  constant123_outs_valid;
  wire  constant123_outs_ready;
  wire [15:0] constant223_outs;
  wire  constant223_outs_valid;
  wire  constant223_outs_ready;
  wire [11:0] constant224_outs;
  wire  constant224_outs_valid;
  wire  constant224_outs_ready;
  wire [11:0] constant126_outs;
  wire  constant126_outs_valid;
  wire  constant126_outs_ready;
  wire [2:0] constant225_outs;
  wire  constant225_outs_valid;
  wire  constant225_outs_ready;
  wire [6:0] constant226_outs;
  wire  constant226_outs_valid;
  wire  constant226_outs_ready;
  wire  source3_outs_valid;
  wire  source3_outs_ready;
  wire [2:0] constant227_outs;
  wire  constant227_outs_valid;
  wire  constant227_outs_ready;
  wire [0:0] cmpi2_result;
  wire  cmpi2_result_valid;
  wire  cmpi2_result_ready;
  wire [0:0] fork9_outs_0;
  wire  fork9_outs_0_valid;
  wire  fork9_outs_0_ready;
  wire [0:0] fork9_outs_1;
  wire  fork9_outs_1_valid;
  wire  fork9_outs_1_ready;
  wire [0:0] fork9_outs_2;
  wire  fork9_outs_2_valid;
  wire  fork9_outs_2_ready;
  wire [0:0] fork9_outs_3;
  wire  fork9_outs_3_valid;
  wire  fork9_outs_3_ready;
  wire [0:0] fork9_outs_4;
  wire  fork9_outs_4_valid;
  wire  fork9_outs_4_ready;
  wire [0:0] fork9_outs_5;
  wire  fork9_outs_5_valid;
  wire  fork9_outs_5_ready;
  wire [0:0] fork9_outs_6;
  wire  fork9_outs_6_valid;
  wire  fork9_outs_6_ready;
  wire [0:0] fork9_outs_7;
  wire  fork9_outs_7_valid;
  wire  fork9_outs_7_ready;
  wire [0:0] fork9_outs_8;
  wire  fork9_outs_8_valid;
  wire  fork9_outs_8_ready;
  wire [0:0] fork9_outs_9;
  wire  fork9_outs_9_valid;
  wire  fork9_outs_9_ready;
  wire [0:0] fork9_outs_10;
  wire  fork9_outs_10_valid;
  wire  fork9_outs_10_ready;
  wire [0:0] fork9_outs_11;
  wire  fork9_outs_11_valid;
  wire  fork9_outs_11_ready;
  wire [0:0] fork9_outs_12;
  wire  fork9_outs_12_valid;
  wire  fork9_outs_12_ready;
  wire [0:0] fork9_outs_13;
  wire  fork9_outs_13_valid;
  wire  fork9_outs_13_ready;
  wire [35:0] cond_br36_trueOut;
  wire  cond_br36_trueOut_valid;
  wire  cond_br36_trueOut_ready;
  wire [35:0] cond_br36_falseOut;
  wire  cond_br36_falseOut_valid;
  wire  cond_br36_falseOut_ready;
  wire [32:0] cond_br37_trueOut;
  wire  cond_br37_trueOut_valid;
  wire  cond_br37_trueOut_ready;
  wire [32:0] cond_br37_falseOut;
  wire  cond_br37_falseOut_valid;
  wire  cond_br37_falseOut_ready;
  wire [33:0] extsi106_outs;
  wire  extsi106_outs_valid;
  wire  extsi106_outs_ready;
  wire [29:0] cond_br38_trueOut;
  wire  cond_br38_trueOut_valid;
  wire  cond_br38_trueOut_ready;
  wire [29:0] cond_br38_falseOut;
  wire  cond_br38_falseOut_valid;
  wire  cond_br38_falseOut_ready;
  wire [25:0] cond_br39_trueOut;
  wire  cond_br39_trueOut_valid;
  wire  cond_br39_trueOut_ready;
  wire [25:0] cond_br39_falseOut;
  wire  cond_br39_falseOut_valid;
  wire  cond_br39_falseOut_ready;
  wire [26:0] extsi107_outs;
  wire  extsi107_outs_valid;
  wire  extsi107_outs_ready;
  wire [21:0] cond_br40_trueOut;
  wire  cond_br40_trueOut_valid;
  wire  cond_br40_trueOut_ready;
  wire [21:0] cond_br40_falseOut;
  wire  cond_br40_falseOut_valid;
  wire  cond_br40_falseOut_ready;
  wire [23:0] extsi108_outs;
  wire  extsi108_outs_valid;
  wire  extsi108_outs_ready;
  wire [20:0] cond_br41_trueOut;
  wire  cond_br41_trueOut_valid;
  wire  cond_br41_trueOut_ready;
  wire [20:0] cond_br41_falseOut;
  wire  cond_br41_falseOut_valid;
  wire  cond_br41_falseOut_ready;
  wire [15:0] cond_br42_trueOut;
  wire  cond_br42_trueOut_valid;
  wire  cond_br42_trueOut_ready;
  wire [15:0] cond_br42_falseOut;
  wire  cond_br42_falseOut_valid;
  wire  cond_br42_falseOut_ready;
  wire [17:0] extsi109_outs;
  wire  extsi109_outs_valid;
  wire  extsi109_outs_ready;
  wire [11:0] cond_br43_trueOut;
  wire  cond_br43_trueOut_valid;
  wire  cond_br43_trueOut_ready;
  wire [11:0] cond_br43_falseOut;
  wire  cond_br43_falseOut_valid;
  wire  cond_br43_falseOut_ready;
  wire [13:0] extsi110_outs;
  wire  extsi110_outs_valid;
  wire  extsi110_outs_ready;
  wire [11:0] cond_br44_trueOut;
  wire  cond_br44_trueOut_valid;
  wire  cond_br44_trueOut_ready;
  wire [11:0] cond_br44_falseOut;
  wire  cond_br44_falseOut_valid;
  wire  cond_br44_falseOut_ready;
  wire [2:0] cond_br45_trueOut;
  wire  cond_br45_trueOut_valid;
  wire  cond_br45_trueOut_ready;
  wire [2:0] cond_br45_falseOut;
  wire  cond_br45_falseOut_valid;
  wire  cond_br45_falseOut_ready;
  wire [7:0] extsi111_outs;
  wire  extsi111_outs_valid;
  wire  extsi111_outs_ready;
  wire [6:0] cond_br46_trueOut;
  wire  cond_br46_trueOut_valid;
  wire  cond_br46_trueOut_ready;
  wire [6:0] cond_br46_falseOut;
  wire  cond_br46_falseOut_valid;
  wire  cond_br46_falseOut_ready;
  wire [7:0] extsi112_outs;
  wire  extsi112_outs_valid;
  wire  extsi112_outs_ready;
  wire [4:0] buffer6_outs;
  wire  buffer6_outs_valid;
  wire  buffer6_outs_ready;
  wire [4:0] buffer7_outs;
  wire  buffer7_outs_valid;
  wire  buffer7_outs_ready;
  wire [4:0] cond_br47_trueOut;
  wire  cond_br47_trueOut_valid;
  wire  cond_br47_trueOut_ready;
  wire [4:0] cond_br47_falseOut;
  wire  cond_br47_falseOut_valid;
  wire  cond_br47_falseOut_ready;
  wire  cond_br48_trueOut_valid;
  wire  cond_br48_trueOut_ready;
  wire  cond_br48_falseOut_valid;
  wire  cond_br48_falseOut_ready;
  wire [2:0] cond_br49_trueOut;
  wire  cond_br49_trueOut_valid;
  wire  cond_br49_trueOut_ready;
  wire [2:0] cond_br49_falseOut;
  wire  cond_br49_falseOut_valid;
  wire  cond_br49_falseOut_ready;
  wire [2:0] buffer14_outs;
  wire  buffer14_outs_valid;
  wire  buffer14_outs_ready;
  wire [2:0] buffer15_outs;
  wire  buffer15_outs_valid;
  wire  buffer15_outs_ready;
  wire [2:0] fork10_outs_0;
  wire  fork10_outs_0_valid;
  wire  fork10_outs_0_ready;
  wire [2:0] fork10_outs_1;
  wire  fork10_outs_1_valid;
  wire  fork10_outs_1_ready;
  wire  buffer16_outs_valid;
  wire  buffer16_outs_ready;
  wire  buffer17_outs_valid;
  wire  buffer17_outs_ready;
  wire  fork11_outs_0_valid;
  wire  fork11_outs_0_ready;
  wire  fork11_outs_1_valid;
  wire  fork11_outs_1_ready;
  wire  fork11_outs_2_valid;
  wire  fork11_outs_2_ready;
  wire  fork11_outs_3_valid;
  wire  fork11_outs_3_ready;
  wire  fork11_outs_4_valid;
  wire  fork11_outs_4_ready;
  wire  fork11_outs_5_valid;
  wire  fork11_outs_5_ready;
  wire  fork11_outs_6_valid;
  wire  fork11_outs_6_ready;
  wire  fork11_outs_7_valid;
  wire  fork11_outs_7_ready;
  wire  fork11_outs_8_valid;
  wire  fork11_outs_8_ready;
  wire  fork11_outs_9_valid;
  wire  fork11_outs_9_ready;
  wire  fork11_outs_10_valid;
  wire  fork11_outs_10_ready;
  wire  fork11_outs_11_valid;
  wire  fork11_outs_11_ready;
  wire [35:0] constant130_outs;
  wire  constant130_outs_valid;
  wire  constant130_outs_ready;
  wire [31:0] constant228_outs;
  wire  constant228_outs_valid;
  wire  constant228_outs_ready;
  wire [29:0] constant132_outs;
  wire  constant132_outs_valid;
  wire  constant132_outs_ready;
  wire [25:0] constant229_outs;
  wire  constant229_outs_valid;
  wire  constant229_outs_ready;
  wire [23:0] constant134_outs;
  wire  constant134_outs_valid;
  wire  constant134_outs_ready;
  wire [20:0] constant135_outs;
  wire  constant135_outs_valid;
  wire  constant135_outs_ready;
  wire [15:0] constant230_outs;
  wire  constant230_outs_valid;
  wire  constant230_outs_ready;
  wire [13:0] constant137_outs;
  wire  constant137_outs_valid;
  wire  constant137_outs_ready;
  wire [11:0] constant138_outs;
  wire  constant138_outs_valid;
  wire  constant138_outs_ready;
  wire [5:0] constant231_outs;
  wire  constant231_outs_valid;
  wire  constant231_outs_ready;
  wire [5:0] constant232_outs;
  wire  constant232_outs_valid;
  wire  constant232_outs_ready;
  wire  source4_outs_valid;
  wire  source4_outs_ready;
  wire [2:0] constant233_outs;
  wire  constant233_outs_valid;
  wire  constant233_outs_ready;
  wire [0:0] cmpi3_result;
  wire  cmpi3_result_valid;
  wire  cmpi3_result_ready;
  wire [0:0] fork12_outs_0;
  wire  fork12_outs_0_valid;
  wire  fork12_outs_0_ready;
  wire [0:0] fork12_outs_1;
  wire  fork12_outs_1_valid;
  wire  fork12_outs_1_ready;
  wire [0:0] fork12_outs_2;
  wire  fork12_outs_2_valid;
  wire  fork12_outs_2_ready;
  wire [0:0] fork12_outs_3;
  wire  fork12_outs_3_valid;
  wire  fork12_outs_3_ready;
  wire [0:0] fork12_outs_4;
  wire  fork12_outs_4_valid;
  wire  fork12_outs_4_ready;
  wire [0:0] fork12_outs_5;
  wire  fork12_outs_5_valid;
  wire  fork12_outs_5_ready;
  wire [0:0] fork12_outs_6;
  wire  fork12_outs_6_valid;
  wire  fork12_outs_6_ready;
  wire [0:0] fork12_outs_7;
  wire  fork12_outs_7_valid;
  wire  fork12_outs_7_ready;
  wire [0:0] fork12_outs_8;
  wire  fork12_outs_8_valid;
  wire  fork12_outs_8_ready;
  wire [0:0] fork12_outs_9;
  wire  fork12_outs_9_valid;
  wire  fork12_outs_9_ready;
  wire [0:0] fork12_outs_10;
  wire  fork12_outs_10_valid;
  wire  fork12_outs_10_ready;
  wire [0:0] fork12_outs_11;
  wire  fork12_outs_11_valid;
  wire  fork12_outs_11_ready;
  wire [0:0] fork12_outs_12;
  wire  fork12_outs_12_valid;
  wire  fork12_outs_12_ready;
  wire [0:0] fork12_outs_13;
  wire  fork12_outs_13_valid;
  wire  fork12_outs_13_ready;
  wire [35:0] cond_br50_trueOut;
  wire  cond_br50_trueOut_valid;
  wire  cond_br50_trueOut_ready;
  wire [35:0] cond_br50_falseOut;
  wire  cond_br50_falseOut_valid;
  wire  cond_br50_falseOut_ready;
  wire [31:0] cond_br51_trueOut;
  wire  cond_br51_trueOut_valid;
  wire  cond_br51_trueOut_ready;
  wire [31:0] cond_br51_falseOut;
  wire  cond_br51_falseOut_valid;
  wire  cond_br51_falseOut_ready;
  wire [33:0] extsi113_outs;
  wire  extsi113_outs_valid;
  wire  extsi113_outs_ready;
  wire [29:0] cond_br52_trueOut;
  wire  cond_br52_trueOut_valid;
  wire  cond_br52_trueOut_ready;
  wire [29:0] cond_br52_falseOut;
  wire  cond_br52_falseOut_valid;
  wire  cond_br52_falseOut_ready;
  wire [25:0] cond_br53_trueOut;
  wire  cond_br53_trueOut_valid;
  wire  cond_br53_trueOut_ready;
  wire [25:0] cond_br53_falseOut;
  wire  cond_br53_falseOut_valid;
  wire  cond_br53_falseOut_ready;
  wire [26:0] extsi114_outs;
  wire  extsi114_outs_valid;
  wire  extsi114_outs_ready;
  wire [23:0] cond_br54_trueOut;
  wire  cond_br54_trueOut_valid;
  wire  cond_br54_trueOut_ready;
  wire [23:0] cond_br54_falseOut;
  wire  cond_br54_falseOut_valid;
  wire  cond_br54_falseOut_ready;
  wire [20:0] cond_br55_trueOut;
  wire  cond_br55_trueOut_valid;
  wire  cond_br55_trueOut_ready;
  wire [20:0] cond_br55_falseOut;
  wire  cond_br55_falseOut_valid;
  wire  cond_br55_falseOut_ready;
  wire [15:0] cond_br56_trueOut;
  wire  cond_br56_trueOut_valid;
  wire  cond_br56_trueOut_ready;
  wire [15:0] cond_br56_falseOut;
  wire  cond_br56_falseOut_valid;
  wire  cond_br56_falseOut_ready;
  wire [17:0] extsi115_outs;
  wire  extsi115_outs_valid;
  wire  extsi115_outs_ready;
  wire [13:0] cond_br57_trueOut;
  wire  cond_br57_trueOut_valid;
  wire  cond_br57_trueOut_ready;
  wire [13:0] cond_br57_falseOut;
  wire  cond_br57_falseOut_valid;
  wire  cond_br57_falseOut_ready;
  wire [11:0] cond_br58_trueOut;
  wire  cond_br58_trueOut_valid;
  wire  cond_br58_trueOut_ready;
  wire [11:0] cond_br58_falseOut;
  wire  cond_br58_falseOut_valid;
  wire  cond_br58_falseOut_ready;
  wire [5:0] cond_br59_trueOut;
  wire  cond_br59_trueOut_valid;
  wire  cond_br59_trueOut_ready;
  wire [5:0] cond_br59_falseOut;
  wire  cond_br59_falseOut_valid;
  wire  cond_br59_falseOut_ready;
  wire [7:0] extsi116_outs;
  wire  extsi116_outs_valid;
  wire  extsi116_outs_ready;
  wire [5:0] cond_br60_trueOut;
  wire  cond_br60_trueOut_valid;
  wire  cond_br60_trueOut_ready;
  wire [5:0] cond_br60_falseOut;
  wire  cond_br60_falseOut_valid;
  wire  cond_br60_falseOut_ready;
  wire [7:0] extsi117_outs;
  wire  extsi117_outs_valid;
  wire  extsi117_outs_ready;
  wire [4:0] buffer12_outs;
  wire  buffer12_outs_valid;
  wire  buffer12_outs_ready;
  wire [4:0] buffer13_outs;
  wire  buffer13_outs_valid;
  wire  buffer13_outs_ready;
  wire [4:0] cond_br61_trueOut;
  wire  cond_br61_trueOut_valid;
  wire  cond_br61_trueOut_ready;
  wire [4:0] cond_br61_falseOut;
  wire  cond_br61_falseOut_valid;
  wire  cond_br61_falseOut_ready;
  wire  cond_br62_trueOut_valid;
  wire  cond_br62_trueOut_ready;
  wire  cond_br62_falseOut_valid;
  wire  cond_br62_falseOut_ready;
  wire [2:0] cond_br63_trueOut;
  wire  cond_br63_trueOut_valid;
  wire  cond_br63_trueOut_ready;
  wire [2:0] cond_br63_falseOut;
  wire  cond_br63_falseOut_valid;
  wire  cond_br63_falseOut_ready;
  wire [2:0] buffer20_outs;
  wire  buffer20_outs_valid;
  wire  buffer20_outs_ready;
  wire [2:0] buffer21_outs;
  wire  buffer21_outs_valid;
  wire  buffer21_outs_ready;
  wire [2:0] fork13_outs_0;
  wire  fork13_outs_0_valid;
  wire  fork13_outs_0_ready;
  wire [2:0] fork13_outs_1;
  wire  fork13_outs_1_valid;
  wire  fork13_outs_1_ready;
  wire [3:0] extsi118_outs;
  wire  extsi118_outs_valid;
  wire  extsi118_outs_ready;
  wire  buffer22_outs_valid;
  wire  buffer22_outs_ready;
  wire  buffer23_outs_valid;
  wire  buffer23_outs_ready;
  wire  fork14_outs_0_valid;
  wire  fork14_outs_0_ready;
  wire  fork14_outs_1_valid;
  wire  fork14_outs_1_ready;
  wire  fork14_outs_2_valid;
  wire  fork14_outs_2_ready;
  wire  fork14_outs_3_valid;
  wire  fork14_outs_3_ready;
  wire  fork14_outs_4_valid;
  wire  fork14_outs_4_ready;
  wire  fork14_outs_5_valid;
  wire  fork14_outs_5_ready;
  wire  fork14_outs_6_valid;
  wire  fork14_outs_6_ready;
  wire  fork14_outs_7_valid;
  wire  fork14_outs_7_ready;
  wire  fork14_outs_8_valid;
  wire  fork14_outs_8_ready;
  wire  fork14_outs_9_valid;
  wire  fork14_outs_9_ready;
  wire  fork14_outs_10_valid;
  wire  fork14_outs_10_ready;
  wire  fork14_outs_11_valid;
  wire  fork14_outs_11_ready;
  wire [2:0] constant234_outs;
  wire  constant234_outs_valid;
  wire  constant234_outs_ready;
  wire [35:0] constant143_outs;
  wire  constant143_outs_valid;
  wire  constant143_outs_ready;
  wire [30:0] constant235_outs;
  wire  constant235_outs_valid;
  wire  constant235_outs_ready;
  wire [29:0] constant145_outs;
  wire  constant145_outs_valid;
  wire  constant145_outs_ready;
  wire [24:0] constant236_outs;
  wire  constant236_outs_valid;
  wire  constant236_outs_ready;
  wire [23:0] constant147_outs;
  wire  constant147_outs_valid;
  wire  constant147_outs_ready;
  wire [15:0] constant237_outs;
  wire  constant237_outs_valid;
  wire  constant237_outs_ready;
  wire [12:0] constant238_outs;
  wire  constant238_outs_valid;
  wire  constant238_outs_ready;
  wire [13:0] constant150_outs;
  wire  constant150_outs_valid;
  wire  constant150_outs_ready;
  wire [11:0] constant151_outs;
  wire  constant151_outs_valid;
  wire  constant151_outs_ready;
  wire [6:0] constant239_outs;
  wire  constant239_outs_valid;
  wire  constant239_outs_ready;
  wire  source5_outs_valid;
  wire  source5_outs_ready;
  wire [3:0] constant240_outs;
  wire  constant240_outs_valid;
  wire  constant240_outs_ready;
  wire [0:0] cmpi4_result;
  wire  cmpi4_result_valid;
  wire  cmpi4_result_ready;
  wire [0:0] fork15_outs_0;
  wire  fork15_outs_0_valid;
  wire  fork15_outs_0_ready;
  wire [0:0] fork15_outs_1;
  wire  fork15_outs_1_valid;
  wire  fork15_outs_1_ready;
  wire [0:0] fork15_outs_2;
  wire  fork15_outs_2_valid;
  wire  fork15_outs_2_ready;
  wire [0:0] fork15_outs_3;
  wire  fork15_outs_3_valid;
  wire  fork15_outs_3_ready;
  wire [0:0] fork15_outs_4;
  wire  fork15_outs_4_valid;
  wire  fork15_outs_4_ready;
  wire [0:0] fork15_outs_5;
  wire  fork15_outs_5_valid;
  wire  fork15_outs_5_ready;
  wire [0:0] fork15_outs_6;
  wire  fork15_outs_6_valid;
  wire  fork15_outs_6_ready;
  wire [0:0] fork15_outs_7;
  wire  fork15_outs_7_valid;
  wire  fork15_outs_7_ready;
  wire [0:0] fork15_outs_8;
  wire  fork15_outs_8_valid;
  wire  fork15_outs_8_ready;
  wire [0:0] fork15_outs_9;
  wire  fork15_outs_9_valid;
  wire  fork15_outs_9_ready;
  wire [0:0] fork15_outs_10;
  wire  fork15_outs_10_valid;
  wire  fork15_outs_10_ready;
  wire [0:0] fork15_outs_11;
  wire  fork15_outs_11_valid;
  wire  fork15_outs_11_ready;
  wire [0:0] fork15_outs_12;
  wire  fork15_outs_12_valid;
  wire  fork15_outs_12_ready;
  wire [0:0] fork15_outs_13;
  wire  fork15_outs_13_valid;
  wire  fork15_outs_13_ready;
  wire [35:0] cond_br64_trueOut;
  wire  cond_br64_trueOut_valid;
  wire  cond_br64_trueOut_ready;
  wire [35:0] cond_br64_falseOut;
  wire  cond_br64_falseOut_valid;
  wire  cond_br64_falseOut_ready;
  wire [30:0] cond_br65_trueOut;
  wire  cond_br65_trueOut_valid;
  wire  cond_br65_trueOut_ready;
  wire [30:0] cond_br65_falseOut;
  wire  cond_br65_falseOut_valid;
  wire  cond_br65_falseOut_ready;
  wire [33:0] extsi119_outs;
  wire  extsi119_outs_valid;
  wire  extsi119_outs_ready;
  wire [29:0] cond_br66_trueOut;
  wire  cond_br66_trueOut_valid;
  wire  cond_br66_trueOut_ready;
  wire [29:0] cond_br66_falseOut;
  wire  cond_br66_falseOut_valid;
  wire  cond_br66_falseOut_ready;
  wire [24:0] cond_br67_trueOut;
  wire  cond_br67_trueOut_valid;
  wire  cond_br67_trueOut_ready;
  wire [24:0] cond_br67_falseOut;
  wire  cond_br67_falseOut_valid;
  wire  cond_br67_falseOut_ready;
  wire [26:0] extsi120_outs;
  wire  extsi120_outs_valid;
  wire  extsi120_outs_ready;
  wire [23:0] cond_br68_trueOut;
  wire  cond_br68_trueOut_valid;
  wire  cond_br68_trueOut_ready;
  wire [23:0] cond_br68_falseOut;
  wire  cond_br68_falseOut_valid;
  wire  cond_br68_falseOut_ready;
  wire [15:0] cond_br69_trueOut;
  wire  cond_br69_trueOut_valid;
  wire  cond_br69_trueOut_ready;
  wire [15:0] cond_br69_falseOut;
  wire  cond_br69_falseOut_valid;
  wire  cond_br69_falseOut_ready;
  wire [20:0] extsi121_outs;
  wire  extsi121_outs_valid;
  wire  extsi121_outs_ready;
  wire [12:0] cond_br70_trueOut;
  wire  cond_br70_trueOut_valid;
  wire  cond_br70_trueOut_ready;
  wire [12:0] cond_br70_falseOut;
  wire  cond_br70_falseOut_valid;
  wire  cond_br70_falseOut_ready;
  wire [17:0] extsi122_outs;
  wire  extsi122_outs_valid;
  wire  extsi122_outs_ready;
  wire [13:0] cond_br71_trueOut;
  wire  cond_br71_trueOut_valid;
  wire  cond_br71_trueOut_ready;
  wire [13:0] cond_br71_falseOut;
  wire  cond_br71_falseOut_valid;
  wire  cond_br71_falseOut_ready;
  wire [11:0] cond_br72_trueOut;
  wire  cond_br72_trueOut_valid;
  wire  cond_br72_trueOut_ready;
  wire [11:0] cond_br72_falseOut;
  wire  cond_br72_falseOut_valid;
  wire  cond_br72_falseOut_ready;
  wire [2:0] cond_br73_trueOut;
  wire  cond_br73_trueOut_valid;
  wire  cond_br73_trueOut_ready;
  wire [2:0] cond_br73_falseOut;
  wire  cond_br73_falseOut_valid;
  wire  cond_br73_falseOut_ready;
  wire [7:0] extsi123_outs;
  wire  extsi123_outs_valid;
  wire  extsi123_outs_ready;
  wire [6:0] cond_br74_trueOut;
  wire  cond_br74_trueOut_valid;
  wire  cond_br74_trueOut_ready;
  wire [6:0] cond_br74_falseOut;
  wire  cond_br74_falseOut_valid;
  wire  cond_br74_falseOut_ready;
  wire [7:0] extsi124_outs;
  wire  extsi124_outs_valid;
  wire  extsi124_outs_ready;
  wire [4:0] buffer18_outs;
  wire  buffer18_outs_valid;
  wire  buffer18_outs_ready;
  wire [4:0] buffer19_outs;
  wire  buffer19_outs_valid;
  wire  buffer19_outs_ready;
  wire [4:0] cond_br75_trueOut;
  wire  cond_br75_trueOut_valid;
  wire  cond_br75_trueOut_ready;
  wire [4:0] cond_br75_falseOut;
  wire  cond_br75_falseOut_valid;
  wire  cond_br75_falseOut_ready;
  wire  cond_br76_trueOut_valid;
  wire  cond_br76_trueOut_ready;
  wire  cond_br76_falseOut_valid;
  wire  cond_br76_falseOut_ready;
  wire [2:0] cond_br77_trueOut;
  wire  cond_br77_trueOut_valid;
  wire  cond_br77_trueOut_ready;
  wire [2:0] cond_br77_falseOut;
  wire  cond_br77_falseOut_valid;
  wire  cond_br77_falseOut_ready;
  wire [2:0] buffer26_outs;
  wire  buffer26_outs_valid;
  wire  buffer26_outs_ready;
  wire [2:0] buffer27_outs;
  wire  buffer27_outs_valid;
  wire  buffer27_outs_ready;
  wire [2:0] fork16_outs_0;
  wire  fork16_outs_0_valid;
  wire  fork16_outs_0_ready;
  wire [2:0] fork16_outs_1;
  wire  fork16_outs_1_valid;
  wire  fork16_outs_1_ready;
  wire [3:0] extsi125_outs;
  wire  extsi125_outs_valid;
  wire  extsi125_outs_ready;
  wire  buffer28_outs_valid;
  wire  buffer28_outs_ready;
  wire  buffer29_outs_valid;
  wire  buffer29_outs_ready;
  wire  fork17_outs_0_valid;
  wire  fork17_outs_0_ready;
  wire  fork17_outs_1_valid;
  wire  fork17_outs_1_ready;
  wire  fork17_outs_2_valid;
  wire  fork17_outs_2_ready;
  wire  fork17_outs_3_valid;
  wire  fork17_outs_3_ready;
  wire  fork17_outs_4_valid;
  wire  fork17_outs_4_ready;
  wire  fork17_outs_5_valid;
  wire  fork17_outs_5_ready;
  wire  fork17_outs_6_valid;
  wire  fork17_outs_6_ready;
  wire  fork17_outs_7_valid;
  wire  fork17_outs_7_ready;
  wire  fork17_outs_8_valid;
  wire  fork17_outs_8_ready;
  wire  fork17_outs_9_valid;
  wire  fork17_outs_9_ready;
  wire  fork17_outs_10_valid;
  wire  fork17_outs_10_ready;
  wire  fork17_outs_11_valid;
  wire  fork17_outs_11_ready;
  wire [7:0] constant154_outs;
  wire  constant154_outs_valid;
  wire  constant154_outs_ready;
  wire [35:0] constant155_outs;
  wire  constant155_outs_valid;
  wire  constant155_outs_ready;
  wire [29:0] constant241_outs;
  wire  constant241_outs_valid;
  wire  constant241_outs_ready;
  wire [29:0] constant157_outs;
  wire  constant157_outs_valid;
  wire  constant157_outs_ready;
  wire [23:0] constant242_outs;
  wire  constant242_outs_valid;
  wire  constant242_outs_ready;
  wire [23:0] constant159_outs;
  wire  constant159_outs_valid;
  wire  constant159_outs_ready;
  wire [16:0] constant243_outs;
  wire  constant243_outs_valid;
  wire  constant243_outs_ready;
  wire [17:0] constant161_outs;
  wire  constant161_outs_valid;
  wire  constant161_outs_ready;
  wire [13:0] constant162_outs;
  wire  constant162_outs_valid;
  wire  constant162_outs_ready;
  wire [8:0] constant244_outs;
  wire  constant244_outs_valid;
  wire  constant244_outs_ready;
  wire [5:0] constant245_outs;
  wire  constant245_outs_valid;
  wire  constant245_outs_ready;
  wire  source6_outs_valid;
  wire  source6_outs_ready;
  wire [3:0] constant246_outs;
  wire  constant246_outs_valid;
  wire  constant246_outs_ready;
  wire [0:0] cmpi5_result;
  wire  cmpi5_result_valid;
  wire  cmpi5_result_ready;
  wire [0:0] fork18_outs_0;
  wire  fork18_outs_0_valid;
  wire  fork18_outs_0_ready;
  wire [0:0] fork18_outs_1;
  wire  fork18_outs_1_valid;
  wire  fork18_outs_1_ready;
  wire [0:0] fork18_outs_2;
  wire  fork18_outs_2_valid;
  wire  fork18_outs_2_ready;
  wire [0:0] fork18_outs_3;
  wire  fork18_outs_3_valid;
  wire  fork18_outs_3_ready;
  wire [0:0] fork18_outs_4;
  wire  fork18_outs_4_valid;
  wire  fork18_outs_4_ready;
  wire [0:0] fork18_outs_5;
  wire  fork18_outs_5_valid;
  wire  fork18_outs_5_ready;
  wire [0:0] fork18_outs_6;
  wire  fork18_outs_6_valid;
  wire  fork18_outs_6_ready;
  wire [0:0] fork18_outs_7;
  wire  fork18_outs_7_valid;
  wire  fork18_outs_7_ready;
  wire [0:0] fork18_outs_8;
  wire  fork18_outs_8_valid;
  wire  fork18_outs_8_ready;
  wire [0:0] fork18_outs_9;
  wire  fork18_outs_9_valid;
  wire  fork18_outs_9_ready;
  wire [0:0] fork18_outs_10;
  wire  fork18_outs_10_valid;
  wire  fork18_outs_10_ready;
  wire [0:0] fork18_outs_11;
  wire  fork18_outs_11_valid;
  wire  fork18_outs_11_ready;
  wire [0:0] fork18_outs_12;
  wire  fork18_outs_12_valid;
  wire  fork18_outs_12_ready;
  wire [0:0] fork18_outs_13;
  wire  fork18_outs_13_valid;
  wire  fork18_outs_13_ready;
  wire [35:0] cond_br78_trueOut;
  wire  cond_br78_trueOut_valid;
  wire  cond_br78_trueOut_ready;
  wire [35:0] cond_br78_falseOut;
  wire  cond_br78_falseOut_valid;
  wire  cond_br78_falseOut_ready;
  wire [29:0] cond_br79_trueOut;
  wire  cond_br79_trueOut_valid;
  wire  cond_br79_trueOut_ready;
  wire [29:0] cond_br79_falseOut;
  wire  cond_br79_falseOut_valid;
  wire  cond_br79_falseOut_ready;
  wire [33:0] extsi126_outs;
  wire  extsi126_outs_valid;
  wire  extsi126_outs_ready;
  wire [29:0] cond_br80_trueOut;
  wire  cond_br80_trueOut_valid;
  wire  cond_br80_trueOut_ready;
  wire [29:0] cond_br80_falseOut;
  wire  cond_br80_falseOut_valid;
  wire  cond_br80_falseOut_ready;
  wire [23:0] cond_br81_trueOut;
  wire  cond_br81_trueOut_valid;
  wire  cond_br81_trueOut_ready;
  wire [23:0] cond_br81_falseOut;
  wire  cond_br81_falseOut_valid;
  wire  cond_br81_falseOut_ready;
  wire [26:0] extsi127_outs;
  wire  extsi127_outs_valid;
  wire  extsi127_outs_ready;
  wire [23:0] cond_br82_trueOut;
  wire  cond_br82_trueOut_valid;
  wire  cond_br82_trueOut_ready;
  wire [23:0] cond_br82_falseOut;
  wire  cond_br82_falseOut_valid;
  wire  cond_br82_falseOut_ready;
  wire [16:0] cond_br83_trueOut;
  wire  cond_br83_trueOut_valid;
  wire  cond_br83_trueOut_ready;
  wire [16:0] cond_br83_falseOut;
  wire  cond_br83_falseOut_valid;
  wire  cond_br83_falseOut_ready;
  wire [20:0] extsi128_outs;
  wire  extsi128_outs_valid;
  wire  extsi128_outs_ready;
  wire [17:0] cond_br84_trueOut;
  wire  cond_br84_trueOut_valid;
  wire  cond_br84_trueOut_ready;
  wire [17:0] cond_br84_falseOut;
  wire  cond_br84_falseOut_valid;
  wire  cond_br84_falseOut_ready;
  wire [13:0] cond_br85_trueOut;
  wire  cond_br85_trueOut_valid;
  wire  cond_br85_trueOut_ready;
  wire [13:0] cond_br85_falseOut;
  wire  cond_br85_falseOut_valid;
  wire  cond_br85_falseOut_ready;
  wire [8:0] cond_br86_trueOut;
  wire  cond_br86_trueOut_valid;
  wire  cond_br86_trueOut_ready;
  wire [8:0] cond_br86_falseOut;
  wire  cond_br86_falseOut_valid;
  wire  cond_br86_falseOut_ready;
  wire [11:0] extsi129_outs;
  wire  extsi129_outs_valid;
  wire  extsi129_outs_ready;
  wire [5:0] cond_br87_trueOut;
  wire  cond_br87_trueOut_valid;
  wire  cond_br87_trueOut_ready;
  wire [5:0] cond_br87_falseOut;
  wire  cond_br87_falseOut_valid;
  wire  cond_br87_falseOut_ready;
  wire [7:0] extsi130_outs;
  wire  extsi130_outs_valid;
  wire  extsi130_outs_ready;
  wire [7:0] cond_br88_trueOut;
  wire  cond_br88_trueOut_valid;
  wire  cond_br88_trueOut_ready;
  wire [7:0] cond_br88_falseOut;
  wire  cond_br88_falseOut_valid;
  wire  cond_br88_falseOut_ready;
  wire [4:0] buffer24_outs;
  wire  buffer24_outs_valid;
  wire  buffer24_outs_ready;
  wire [4:0] buffer25_outs;
  wire  buffer25_outs_valid;
  wire  buffer25_outs_ready;
  wire [4:0] cond_br89_trueOut;
  wire  cond_br89_trueOut_valid;
  wire  cond_br89_trueOut_ready;
  wire [4:0] cond_br89_falseOut;
  wire  cond_br89_falseOut_valid;
  wire  cond_br89_falseOut_ready;
  wire  cond_br90_trueOut_valid;
  wire  cond_br90_trueOut_ready;
  wire  cond_br90_falseOut_valid;
  wire  cond_br90_falseOut_ready;
  wire [2:0] cond_br91_trueOut;
  wire  cond_br91_trueOut_valid;
  wire  cond_br91_trueOut_ready;
  wire [2:0] cond_br91_falseOut;
  wire  cond_br91_falseOut_valid;
  wire  cond_br91_falseOut_ready;
  wire [2:0] buffer32_outs;
  wire  buffer32_outs_valid;
  wire  buffer32_outs_ready;
  wire [2:0] buffer33_outs;
  wire  buffer33_outs_valid;
  wire  buffer33_outs_ready;
  wire [2:0] fork19_outs_0;
  wire  fork19_outs_0_valid;
  wire  fork19_outs_0_ready;
  wire [2:0] fork19_outs_1;
  wire  fork19_outs_1_valid;
  wire  fork19_outs_1_ready;
  wire [3:0] extsi131_outs;
  wire  extsi131_outs_valid;
  wire  extsi131_outs_ready;
  wire  buffer34_outs_valid;
  wire  buffer34_outs_ready;
  wire  buffer35_outs_valid;
  wire  buffer35_outs_ready;
  wire  fork20_outs_0_valid;
  wire  fork20_outs_0_ready;
  wire  fork20_outs_1_valid;
  wire  fork20_outs_1_ready;
  wire  fork20_outs_2_valid;
  wire  fork20_outs_2_ready;
  wire  fork20_outs_3_valid;
  wire  fork20_outs_3_ready;
  wire  fork20_outs_4_valid;
  wire  fork20_outs_4_ready;
  wire  fork20_outs_5_valid;
  wire  fork20_outs_5_ready;
  wire  fork20_outs_6_valid;
  wire  fork20_outs_6_ready;
  wire  fork20_outs_7_valid;
  wire  fork20_outs_7_ready;
  wire  fork20_outs_8_valid;
  wire  fork20_outs_8_ready;
  wire  fork20_outs_9_valid;
  wire  fork20_outs_9_ready;
  wire  fork20_outs_10_valid;
  wire  fork20_outs_10_ready;
  wire  fork20_outs_11_valid;
  wire  fork20_outs_11_ready;
  wire [35:0] constant166_outs;
  wire  constant166_outs_valid;
  wire  constant166_outs_ready;
  wire [28:0] constant247_outs;
  wire  constant247_outs_valid;
  wire  constant247_outs_ready;
  wire [29:0] constant168_outs;
  wire  constant168_outs_valid;
  wire  constant168_outs_ready;
  wire [22:0] constant248_outs;
  wire  constant248_outs_valid;
  wire  constant248_outs_ready;
  wire [23:0] constant170_outs;
  wire  constant170_outs_valid;
  wire  constant170_outs_ready;
  wire [15:0] constant249_outs;
  wire  constant249_outs_valid;
  wire  constant249_outs_ready;
  wire [17:0] constant172_outs;
  wire  constant172_outs_valid;
  wire  constant172_outs_ready;
  wire [5:0] constant250_outs;
  wire  constant250_outs_valid;
  wire  constant250_outs_ready;
  wire [11:0] constant174_outs;
  wire  constant174_outs_valid;
  wire  constant174_outs_ready;
  wire [7:0] constant175_outs;
  wire  constant175_outs_valid;
  wire  constant175_outs_ready;
  wire [4:0] constant251_outs;
  wire  constant251_outs_valid;
  wire  constant251_outs_ready;
  wire  source7_outs_valid;
  wire  source7_outs_ready;
  wire [3:0] constant252_outs;
  wire  constant252_outs_valid;
  wire  constant252_outs_ready;
  wire [0:0] cmpi6_result;
  wire  cmpi6_result_valid;
  wire  cmpi6_result_ready;
  wire [0:0] fork21_outs_0;
  wire  fork21_outs_0_valid;
  wire  fork21_outs_0_ready;
  wire [0:0] fork21_outs_1;
  wire  fork21_outs_1_valid;
  wire  fork21_outs_1_ready;
  wire [0:0] fork21_outs_2;
  wire  fork21_outs_2_valid;
  wire  fork21_outs_2_ready;
  wire [0:0] fork21_outs_3;
  wire  fork21_outs_3_valid;
  wire  fork21_outs_3_ready;
  wire [0:0] fork21_outs_4;
  wire  fork21_outs_4_valid;
  wire  fork21_outs_4_ready;
  wire [0:0] fork21_outs_5;
  wire  fork21_outs_5_valid;
  wire  fork21_outs_5_ready;
  wire [0:0] fork21_outs_6;
  wire  fork21_outs_6_valid;
  wire  fork21_outs_6_ready;
  wire [0:0] fork21_outs_7;
  wire  fork21_outs_7_valid;
  wire  fork21_outs_7_ready;
  wire [0:0] fork21_outs_8;
  wire  fork21_outs_8_valid;
  wire  fork21_outs_8_ready;
  wire [0:0] fork21_outs_9;
  wire  fork21_outs_9_valid;
  wire  fork21_outs_9_ready;
  wire [0:0] fork21_outs_10;
  wire  fork21_outs_10_valid;
  wire  fork21_outs_10_ready;
  wire [0:0] fork21_outs_11;
  wire  fork21_outs_11_valid;
  wire  fork21_outs_11_ready;
  wire [0:0] fork21_outs_12;
  wire  fork21_outs_12_valid;
  wire  fork21_outs_12_ready;
  wire [0:0] fork21_outs_13;
  wire  fork21_outs_13_valid;
  wire  fork21_outs_13_ready;
  wire [35:0] cond_br92_trueOut;
  wire  cond_br92_trueOut_valid;
  wire  cond_br92_trueOut_ready;
  wire [35:0] cond_br92_falseOut;
  wire  cond_br92_falseOut_valid;
  wire  cond_br92_falseOut_ready;
  wire [28:0] cond_br93_trueOut;
  wire  cond_br93_trueOut_valid;
  wire  cond_br93_trueOut_ready;
  wire [28:0] cond_br93_falseOut;
  wire  cond_br93_falseOut_valid;
  wire  cond_br93_falseOut_ready;
  wire [33:0] extsi132_outs;
  wire  extsi132_outs_valid;
  wire  extsi132_outs_ready;
  wire [29:0] cond_br94_trueOut;
  wire  cond_br94_trueOut_valid;
  wire  cond_br94_trueOut_ready;
  wire [29:0] cond_br94_falseOut;
  wire  cond_br94_falseOut_valid;
  wire  cond_br94_falseOut_ready;
  wire [22:0] cond_br95_trueOut;
  wire  cond_br95_trueOut_valid;
  wire  cond_br95_trueOut_ready;
  wire [22:0] cond_br95_falseOut;
  wire  cond_br95_falseOut_valid;
  wire  cond_br95_falseOut_ready;
  wire [26:0] extsi133_outs;
  wire  extsi133_outs_valid;
  wire  extsi133_outs_ready;
  wire [23:0] cond_br96_trueOut;
  wire  cond_br96_trueOut_valid;
  wire  cond_br96_trueOut_ready;
  wire [23:0] cond_br96_falseOut;
  wire  cond_br96_falseOut_valid;
  wire  cond_br96_falseOut_ready;
  wire [15:0] cond_br97_trueOut;
  wire  cond_br97_trueOut_valid;
  wire  cond_br97_trueOut_ready;
  wire [15:0] cond_br97_falseOut;
  wire  cond_br97_falseOut_valid;
  wire  cond_br97_falseOut_ready;
  wire [20:0] extsi134_outs;
  wire  extsi134_outs_valid;
  wire  extsi134_outs_ready;
  wire [17:0] cond_br98_trueOut;
  wire  cond_br98_trueOut_valid;
  wire  cond_br98_trueOut_ready;
  wire [17:0] cond_br98_falseOut;
  wire  cond_br98_falseOut_valid;
  wire  cond_br98_falseOut_ready;
  wire [5:0] cond_br99_trueOut;
  wire  cond_br99_trueOut_valid;
  wire  cond_br99_trueOut_ready;
  wire [5:0] cond_br99_falseOut;
  wire  cond_br99_falseOut_valid;
  wire  cond_br99_falseOut_ready;
  wire [13:0] extsi135_outs;
  wire  extsi135_outs_valid;
  wire  extsi135_outs_ready;
  wire [11:0] cond_br100_trueOut;
  wire  cond_br100_trueOut_valid;
  wire  cond_br100_trueOut_ready;
  wire [11:0] cond_br100_falseOut;
  wire  cond_br100_falseOut_valid;
  wire  cond_br100_falseOut_ready;
  wire [7:0] cond_br101_trueOut;
  wire  cond_br101_trueOut_valid;
  wire  cond_br101_trueOut_ready;
  wire [7:0] cond_br101_falseOut;
  wire  cond_br101_falseOut_valid;
  wire  cond_br101_falseOut_ready;
  wire [4:0] cond_br102_trueOut;
  wire  cond_br102_trueOut_valid;
  wire  cond_br102_trueOut_ready;
  wire [4:0] cond_br102_falseOut;
  wire  cond_br102_falseOut_valid;
  wire  cond_br102_falseOut_ready;
  wire [7:0] extsi136_outs;
  wire  extsi136_outs_valid;
  wire  extsi136_outs_ready;
  wire [4:0] buffer30_outs;
  wire  buffer30_outs_valid;
  wire  buffer30_outs_ready;
  wire [4:0] buffer31_outs;
  wire  buffer31_outs_valid;
  wire  buffer31_outs_ready;
  wire [4:0] cond_br103_trueOut;
  wire  cond_br103_trueOut_valid;
  wire  cond_br103_trueOut_ready;
  wire [4:0] cond_br103_falseOut;
  wire  cond_br103_falseOut_valid;
  wire  cond_br103_falseOut_ready;
  wire  cond_br104_trueOut_valid;
  wire  cond_br104_trueOut_ready;
  wire  cond_br104_falseOut_valid;
  wire  cond_br104_falseOut_ready;
  wire [2:0] cond_br105_trueOut;
  wire  cond_br105_trueOut_valid;
  wire  cond_br105_trueOut_ready;
  wire [2:0] cond_br105_falseOut;
  wire  cond_br105_falseOut_valid;
  wire  cond_br105_falseOut_ready;
  wire [2:0] buffer38_outs;
  wire  buffer38_outs_valid;
  wire  buffer38_outs_ready;
  wire [2:0] buffer39_outs;
  wire  buffer39_outs_valid;
  wire  buffer39_outs_ready;
  wire [3:0] extsi137_outs;
  wire  extsi137_outs_valid;
  wire  extsi137_outs_ready;
  wire  buffer40_outs_valid;
  wire  buffer40_outs_ready;
  wire  buffer41_outs_valid;
  wire  buffer41_outs_ready;
  wire  fork22_outs_0_valid;
  wire  fork22_outs_0_ready;
  wire  fork22_outs_1_valid;
  wire  fork22_outs_1_ready;
  wire  fork22_outs_2_valid;
  wire  fork22_outs_2_ready;
  wire  fork22_outs_3_valid;
  wire  fork22_outs_3_ready;
  wire  fork22_outs_4_valid;
  wire  fork22_outs_4_ready;
  wire  fork22_outs_5_valid;
  wire  fork22_outs_5_ready;
  wire  fork22_outs_6_valid;
  wire  fork22_outs_6_ready;
  wire  fork22_outs_7_valid;
  wire  fork22_outs_7_ready;
  wire  fork22_outs_8_valid;
  wire  fork22_outs_8_ready;
  wire  fork22_outs_9_valid;
  wire  fork22_outs_9_ready;
  wire  fork22_outs_10_valid;
  wire  fork22_outs_10_ready;
  wire  fork22_outs_11_valid;
  wire  fork22_outs_11_ready;
  wire  fork22_outs_12_valid;
  wire  fork22_outs_12_ready;
  wire  fork22_outs_13_valid;
  wire  fork22_outs_13_ready;
  wire  fork22_outs_14_valid;
  wire  fork22_outs_14_ready;
  wire  fork22_outs_15_valid;
  wire  fork22_outs_15_ready;
  wire  fork22_outs_16_valid;
  wire  fork22_outs_16_ready;
  wire  fork22_outs_17_valid;
  wire  fork22_outs_17_ready;
  wire  fork22_outs_18_valid;
  wire  fork22_outs_18_ready;
  wire  fork22_outs_19_valid;
  wire  fork22_outs_19_ready;
  wire  fork22_outs_20_valid;
  wire  fork22_outs_20_ready;
  wire  fork22_outs_21_valid;
  wire  fork22_outs_21_ready;
  wire  fork22_outs_22_valid;
  wire  fork22_outs_22_ready;
  wire [33:0] constant253_outs;
  wire  constant253_outs_valid;
  wire  constant253_outs_ready;
  wire [33:0] constant179_outs;
  wire  constant179_outs_valid;
  wire  constant179_outs_ready;
  wire [29:0] constant180_outs;
  wire  constant180_outs_valid;
  wire  constant180_outs_ready;
  wire [26:0] constant181_outs;
  wire  constant181_outs_valid;
  wire  constant181_outs_ready;
  wire [23:0] constant182_outs;
  wire  constant182_outs_valid;
  wire  constant182_outs_ready;
  wire [20:0] constant183_outs;
  wire  constant183_outs_valid;
  wire  constant183_outs_ready;
  wire [17:0] constant184_outs;
  wire  constant184_outs_valid;
  wire  constant184_outs_ready;
  wire [13:0] constant185_outs;
  wire  constant185_outs_valid;
  wire  constant185_outs_ready;
  wire [11:0] constant186_outs;
  wire  constant186_outs_valid;
  wire  constant186_outs_ready;
  wire [6:0] constant254_outs;
  wire  constant254_outs_valid;
  wire  constant254_outs_ready;
  wire [7:0] constant188_outs;
  wire  constant188_outs_valid;
  wire  constant188_outs_ready;
  wire [35:0] constant189_outs;
  wire  constant189_outs_valid;
  wire  constant189_outs_ready;
  wire [27:0] constant255_outs;
  wire  constant255_outs_valid;
  wire  constant255_outs_ready;
  wire [29:0] constant191_outs;
  wire  constant191_outs_valid;
  wire  constant191_outs_ready;
  wire [21:0] constant256_outs;
  wire  constant256_outs_valid;
  wire  constant256_outs_ready;
  wire [23:0] constant193_outs;
  wire  constant193_outs_valid;
  wire  constant193_outs_ready;
  wire [14:0] constant257_outs;
  wire  constant257_outs_valid;
  wire  constant257_outs_ready;
  wire [17:0] constant195_outs;
  wire  constant195_outs_valid;
  wire  constant195_outs_ready;
  wire [7:0] constant258_outs;
  wire  constant258_outs_valid;
  wire  constant258_outs_ready;
  wire [11:0] constant197_outs;
  wire  constant197_outs_valid;
  wire  constant197_outs_ready;
  wire [7:0] constant198_outs;
  wire  constant198_outs_valid;
  wire  constant198_outs_ready;
  wire [7:0] constant199_outs;
  wire  constant199_outs_valid;
  wire  constant199_outs_ready;
  wire  source8_outs_valid;
  wire  source8_outs_ready;
  wire [3:0] constant259_outs;
  wire  constant259_outs_valid;
  wire  constant259_outs_ready;
  wire [0:0] cmpi7_result;
  wire  cmpi7_result_valid;
  wire  cmpi7_result_ready;
  wire [0:0] fork23_outs_0;
  wire  fork23_outs_0_valid;
  wire  fork23_outs_0_ready;
  wire [0:0] fork23_outs_1;
  wire  fork23_outs_1_valid;
  wire  fork23_outs_1_ready;
  wire [0:0] fork23_outs_2;
  wire  fork23_outs_2_valid;
  wire  fork23_outs_2_ready;
  wire [0:0] fork23_outs_3;
  wire  fork23_outs_3_valid;
  wire  fork23_outs_3_ready;
  wire [0:0] fork23_outs_4;
  wire  fork23_outs_4_valid;
  wire  fork23_outs_4_ready;
  wire [0:0] fork23_outs_5;
  wire  fork23_outs_5_valid;
  wire  fork23_outs_5_ready;
  wire [0:0] fork23_outs_6;
  wire  fork23_outs_6_valid;
  wire  fork23_outs_6_ready;
  wire [0:0] fork23_outs_7;
  wire  fork23_outs_7_valid;
  wire  fork23_outs_7_ready;
  wire [0:0] fork23_outs_8;
  wire  fork23_outs_8_valid;
  wire  fork23_outs_8_ready;
  wire [0:0] fork23_outs_9;
  wire  fork23_outs_9_valid;
  wire  fork23_outs_9_ready;
  wire [0:0] fork23_outs_10;
  wire  fork23_outs_10_valid;
  wire  fork23_outs_10_ready;
  wire [0:0] fork23_outs_11;
  wire  fork23_outs_11_valid;
  wire  fork23_outs_11_ready;
  wire [0:0] fork23_outs_12;
  wire  fork23_outs_12_valid;
  wire  fork23_outs_12_ready;
  wire [0:0] fork23_outs_13;
  wire  fork23_outs_13_valid;
  wire  fork23_outs_13_ready;
  wire [0:0] fork23_outs_14;
  wire  fork23_outs_14_valid;
  wire  fork23_outs_14_ready;
  wire [0:0] fork23_outs_15;
  wire  fork23_outs_15_valid;
  wire  fork23_outs_15_ready;
  wire [0:0] fork23_outs_16;
  wire  fork23_outs_16_valid;
  wire  fork23_outs_16_ready;
  wire [0:0] fork23_outs_17;
  wire  fork23_outs_17_valid;
  wire  fork23_outs_17_ready;
  wire [0:0] fork23_outs_18;
  wire  fork23_outs_18_valid;
  wire  fork23_outs_18_ready;
  wire [0:0] fork23_outs_19;
  wire  fork23_outs_19_valid;
  wire  fork23_outs_19_ready;
  wire [0:0] fork23_outs_20;
  wire  fork23_outs_20_valid;
  wire  fork23_outs_20_ready;
  wire [0:0] fork23_outs_21;
  wire  fork23_outs_21_valid;
  wire  fork23_outs_21_ready;
  wire [0:0] fork23_outs_22;
  wire  fork23_outs_22_valid;
  wire  fork23_outs_22_ready;
  wire [0:0] fork23_outs_23;
  wire  fork23_outs_23_valid;
  wire  fork23_outs_23_ready;
  wire [35:0] cond_br106_trueOut;
  wire  cond_br106_trueOut_valid;
  wire  cond_br106_trueOut_ready;
  wire [35:0] cond_br106_falseOut;
  wire  cond_br106_falseOut_valid;
  wire  cond_br106_falseOut_ready;
  wire [27:0] cond_br107_trueOut;
  wire  cond_br107_trueOut_valid;
  wire  cond_br107_trueOut_ready;
  wire [27:0] cond_br107_falseOut;
  wire  cond_br107_falseOut_valid;
  wire  cond_br107_falseOut_ready;
  wire [33:0] extsi138_outs;
  wire  extsi138_outs_valid;
  wire  extsi138_outs_ready;
  wire [29:0] cond_br108_trueOut;
  wire  cond_br108_trueOut_valid;
  wire  cond_br108_trueOut_ready;
  wire [29:0] cond_br108_falseOut;
  wire  cond_br108_falseOut_valid;
  wire  cond_br108_falseOut_ready;
  wire [21:0] cond_br109_trueOut;
  wire  cond_br109_trueOut_valid;
  wire  cond_br109_trueOut_ready;
  wire [21:0] cond_br109_falseOut;
  wire  cond_br109_falseOut_valid;
  wire  cond_br109_falseOut_ready;
  wire [26:0] extsi139_outs;
  wire  extsi139_outs_valid;
  wire  extsi139_outs_ready;
  wire [23:0] cond_br110_trueOut;
  wire  cond_br110_trueOut_valid;
  wire  cond_br110_trueOut_ready;
  wire [23:0] cond_br110_falseOut;
  wire  cond_br110_falseOut_valid;
  wire  cond_br110_falseOut_ready;
  wire [14:0] cond_br111_trueOut;
  wire  cond_br111_trueOut_valid;
  wire  cond_br111_trueOut_ready;
  wire [14:0] cond_br111_falseOut;
  wire  cond_br111_falseOut_valid;
  wire  cond_br111_falseOut_ready;
  wire [20:0] extsi140_outs;
  wire  extsi140_outs_valid;
  wire  extsi140_outs_ready;
  wire [17:0] cond_br112_trueOut;
  wire  cond_br112_trueOut_valid;
  wire  cond_br112_trueOut_ready;
  wire [17:0] cond_br112_falseOut;
  wire  cond_br112_falseOut_valid;
  wire  cond_br112_falseOut_ready;
  wire [7:0] cond_br113_trueOut;
  wire  cond_br113_trueOut_valid;
  wire  cond_br113_trueOut_ready;
  wire [7:0] cond_br113_falseOut;
  wire  cond_br113_falseOut_valid;
  wire  cond_br113_falseOut_ready;
  wire [13:0] extsi141_outs;
  wire  extsi141_outs_valid;
  wire  extsi141_outs_ready;
  wire [11:0] cond_br114_trueOut;
  wire  cond_br114_trueOut_valid;
  wire  cond_br114_trueOut_ready;
  wire [11:0] cond_br114_falseOut;
  wire  cond_br114_falseOut_valid;
  wire  cond_br114_falseOut_ready;
  wire [7:0] cond_br115_trueOut;
  wire  cond_br115_trueOut_valid;
  wire  cond_br115_trueOut_ready;
  wire [7:0] cond_br115_falseOut;
  wire  cond_br115_falseOut_valid;
  wire  cond_br115_falseOut_ready;
  wire [7:0] cond_br116_trueOut;
  wire  cond_br116_trueOut_valid;
  wire  cond_br116_trueOut_ready;
  wire [7:0] cond_br116_falseOut;
  wire  cond_br116_falseOut_valid;
  wire  cond_br116_falseOut_ready;
  wire [4:0] buffer36_outs;
  wire  buffer36_outs_valid;
  wire  buffer36_outs_ready;
  wire [4:0] buffer37_outs;
  wire  buffer37_outs_valid;
  wire  buffer37_outs_ready;
  wire [4:0] cond_br117_trueOut;
  wire  cond_br117_trueOut_valid;
  wire  cond_br117_trueOut_ready;
  wire [4:0] cond_br117_falseOut;
  wire  cond_br117_falseOut_valid;
  wire  cond_br117_falseOut_ready;
  wire [4:0] fork24_outs_0;
  wire  fork24_outs_0_valid;
  wire  fork24_outs_0_ready;
  wire [4:0] fork24_outs_1;
  wire  fork24_outs_1_valid;
  wire  fork24_outs_1_ready;
  wire  cond_br118_trueOut_valid;
  wire  cond_br118_trueOut_ready;
  wire  cond_br118_falseOut_valid;
  wire  cond_br118_falseOut_ready;
  wire  fork25_outs_0_valid;
  wire  fork25_outs_0_ready;
  wire  fork25_outs_1_valid;
  wire  fork25_outs_1_ready;
  wire [33:0] cond_br119_trueOut;
  wire  cond_br119_trueOut_valid;
  wire  cond_br119_trueOut_ready;
  wire [33:0] cond_br119_falseOut;
  wire  cond_br119_falseOut_valid;
  wire  cond_br119_falseOut_ready;
  wire [35:0] extsi142_outs;
  wire  extsi142_outs_valid;
  wire  extsi142_outs_ready;
  wire [33:0] cond_br120_trueOut;
  wire  cond_br120_trueOut_valid;
  wire  cond_br120_trueOut_ready;
  wire [33:0] cond_br120_falseOut;
  wire  cond_br120_falseOut_valid;
  wire  cond_br120_falseOut_ready;
  wire [29:0] cond_br121_trueOut;
  wire  cond_br121_trueOut_valid;
  wire  cond_br121_trueOut_ready;
  wire [29:0] cond_br121_falseOut;
  wire  cond_br121_falseOut_valid;
  wire  cond_br121_falseOut_ready;
  wire [26:0] cond_br122_trueOut;
  wire  cond_br122_trueOut_valid;
  wire  cond_br122_trueOut_ready;
  wire [26:0] cond_br122_falseOut;
  wire  cond_br122_falseOut_valid;
  wire  cond_br122_falseOut_ready;
  wire [23:0] cond_br123_trueOut;
  wire  cond_br123_trueOut_valid;
  wire  cond_br123_trueOut_ready;
  wire [23:0] cond_br123_falseOut;
  wire  cond_br123_falseOut_valid;
  wire  cond_br123_falseOut_ready;
  wire [20:0] cond_br124_trueOut;
  wire  cond_br124_trueOut_valid;
  wire  cond_br124_trueOut_ready;
  wire [20:0] cond_br124_falseOut;
  wire  cond_br124_falseOut_valid;
  wire  cond_br124_falseOut_ready;
  wire [17:0] cond_br125_trueOut;
  wire  cond_br125_trueOut_valid;
  wire  cond_br125_trueOut_ready;
  wire [17:0] cond_br125_falseOut;
  wire  cond_br125_falseOut_valid;
  wire  cond_br125_falseOut_ready;
  wire [13:0] cond_br126_trueOut;
  wire  cond_br126_trueOut_valid;
  wire  cond_br126_trueOut_ready;
  wire [13:0] cond_br126_falseOut;
  wire  cond_br126_falseOut_valid;
  wire  cond_br126_falseOut_ready;
  wire [11:0] cond_br127_trueOut;
  wire  cond_br127_trueOut_valid;
  wire  cond_br127_trueOut_ready;
  wire [11:0] cond_br127_falseOut;
  wire  cond_br127_falseOut_valid;
  wire  cond_br127_falseOut_ready;
  wire [6:0] cond_br128_trueOut;
  wire  cond_br128_trueOut_valid;
  wire  cond_br128_trueOut_ready;
  wire [6:0] cond_br128_falseOut;
  wire  cond_br128_falseOut_valid;
  wire  cond_br128_falseOut_ready;
  wire [7:0] extsi143_outs;
  wire  extsi143_outs_valid;
  wire  extsi143_outs_ready;
  wire [7:0] cond_br129_trueOut;
  wire  cond_br129_trueOut_valid;
  wire  cond_br129_trueOut_ready;
  wire [7:0] cond_br129_falseOut;
  wire  cond_br129_falseOut_valid;
  wire  cond_br129_falseOut_ready;
  wire [35:0] mux0_outs;
  wire  mux0_outs_valid;
  wire  mux0_outs_ready;
  wire [33:0] mux1_outs;
  wire  mux1_outs_valid;
  wire  mux1_outs_ready;
  wire [29:0] mux2_outs;
  wire  mux2_outs_valid;
  wire  mux2_outs_ready;
  wire [26:0] mux3_outs;
  wire  mux3_outs_valid;
  wire  mux3_outs_ready;
  wire [23:0] mux4_outs;
  wire  mux4_outs_valid;
  wire  mux4_outs_ready;
  wire [20:0] mux5_outs;
  wire  mux5_outs_valid;
  wire  mux5_outs_ready;
  wire [17:0] mux6_outs;
  wire  mux6_outs_valid;
  wire  mux6_outs_ready;
  wire [13:0] mux7_outs;
  wire  mux7_outs_valid;
  wire  mux7_outs_ready;
  wire [11:0] mux8_outs;
  wire  mux8_outs_valid;
  wire  mux8_outs_ready;
  wire [7:0] mux9_outs;
  wire  mux9_outs_valid;
  wire  mux9_outs_ready;
  wire [7:0] mux10_outs;
  wire  mux10_outs_valid;
  wire  mux10_outs_ready;
  wire [7:0] buffer62_outs;
  wire  buffer62_outs_valid;
  wire  buffer62_outs_ready;
  wire [7:0] buffer63_outs;
  wire  buffer63_outs_valid;
  wire  buffer63_outs_ready;
  wire [12:0] extsi144_outs;
  wire  extsi144_outs_valid;
  wire  extsi144_outs_ready;
  wire [4:0] mux11_outs;
  wire  mux11_outs_valid;
  wire  mux11_outs_ready;
  wire [4:0] buffer64_outs;
  wire  buffer64_outs_valid;
  wire  buffer64_outs_ready;
  wire [4:0] buffer65_outs;
  wire  buffer65_outs_valid;
  wire  buffer65_outs_ready;
  wire [4:0] fork26_outs_0;
  wire  fork26_outs_0_valid;
  wire  fork26_outs_0_ready;
  wire [4:0] fork26_outs_1;
  wire  fork26_outs_1_valid;
  wire  fork26_outs_1_ready;
  wire [4:0] fork26_outs_2;
  wire  fork26_outs_2_valid;
  wire  fork26_outs_2_ready;
  wire [4:0] fork26_outs_3;
  wire  fork26_outs_3_valid;
  wire  fork26_outs_3_ready;
  wire [4:0] fork26_outs_4;
  wire  fork26_outs_4_valid;
  wire  fork26_outs_4_ready;
  wire [4:0] fork26_outs_5;
  wire  fork26_outs_5_valid;
  wire  fork26_outs_5_ready;
  wire [4:0] fork26_outs_6;
  wire  fork26_outs_6_valid;
  wire  fork26_outs_6_ready;
  wire [4:0] fork26_outs_7;
  wire  fork26_outs_7_valid;
  wire  fork26_outs_7_ready;
  wire [4:0] fork26_outs_8;
  wire  fork26_outs_8_valid;
  wire  fork26_outs_8_ready;
  wire [4:0] fork26_outs_9;
  wire  fork26_outs_9_valid;
  wire  fork26_outs_9_ready;
  wire  control_merge7_outs_valid;
  wire  control_merge7_outs_ready;
  wire [3:0] control_merge7_index;
  wire  control_merge7_index_valid;
  wire  control_merge7_index_ready;
  wire [3:0] fork27_outs_0;
  wire  fork27_outs_0_valid;
  wire  fork27_outs_0_ready;
  wire [3:0] fork27_outs_1;
  wire  fork27_outs_1_valid;
  wire  fork27_outs_1_ready;
  wire [3:0] fork27_outs_2;
  wire  fork27_outs_2_valid;
  wire  fork27_outs_2_ready;
  wire [3:0] fork27_outs_3;
  wire  fork27_outs_3_valid;
  wire  fork27_outs_3_ready;
  wire [3:0] fork27_outs_4;
  wire  fork27_outs_4_valid;
  wire  fork27_outs_4_ready;
  wire [3:0] fork27_outs_5;
  wire  fork27_outs_5_valid;
  wire  fork27_outs_5_ready;
  wire [3:0] fork27_outs_6;
  wire  fork27_outs_6_valid;
  wire  fork27_outs_6_ready;
  wire [3:0] fork27_outs_7;
  wire  fork27_outs_7_valid;
  wire  fork27_outs_7_ready;
  wire [3:0] fork27_outs_8;
  wire  fork27_outs_8_valid;
  wire  fork27_outs_8_ready;
  wire [3:0] fork27_outs_9;
  wire  fork27_outs_9_valid;
  wire  fork27_outs_9_ready;
  wire [3:0] fork27_outs_10;
  wire  fork27_outs_10_valid;
  wire  fork27_outs_10_ready;
  wire [3:0] fork27_outs_11;
  wire  fork27_outs_11_valid;
  wire  fork27_outs_11_ready;
  wire  buffer66_outs_valid;
  wire  buffer66_outs_ready;
  wire  buffer67_outs_valid;
  wire  buffer67_outs_ready;
  wire  source9_outs_valid;
  wire  source9_outs_ready;
  wire [2:0] constant260_outs;
  wire  constant260_outs_valid;
  wire  constant260_outs_ready;
  wire [2:0] fork28_outs_0;
  wire  fork28_outs_0_valid;
  wire  fork28_outs_0_ready;
  wire [2:0] fork28_outs_1;
  wire  fork28_outs_1_valid;
  wire  fork28_outs_1_ready;
  wire [2:0] fork28_outs_2;
  wire  fork28_outs_2_valid;
  wire  fork28_outs_2_ready;
  wire [2:0] fork28_outs_3;
  wire  fork28_outs_3_valid;
  wire  fork28_outs_3_ready;
  wire [2:0] fork28_outs_4;
  wire  fork28_outs_4_valid;
  wire  fork28_outs_4_ready;
  wire [2:0] fork28_outs_5;
  wire  fork28_outs_5_valid;
  wire  fork28_outs_5_ready;
  wire [2:0] fork28_outs_6;
  wire  fork28_outs_6_valid;
  wire  fork28_outs_6_ready;
  wire [2:0] fork28_outs_7;
  wire  fork28_outs_7_valid;
  wire  fork28_outs_7_ready;
  wire [2:0] fork28_outs_8;
  wire  fork28_outs_8_valid;
  wire  fork28_outs_8_ready;
  wire [2:0] fork28_outs_9;
  wire  fork28_outs_9_valid;
  wire  fork28_outs_9_ready;
  wire [39:0] extsi88_outs;
  wire  extsi88_outs_valid;
  wire  extsi88_outs_ready;
  wire [37:0] extsi89_outs;
  wire  extsi89_outs_valid;
  wire  extsi89_outs_ready;
  wire [33:0] extsi90_outs;
  wire  extsi90_outs_valid;
  wire  extsi90_outs_ready;
  wire [30:0] extsi91_outs;
  wire  extsi91_outs_valid;
  wire  extsi91_outs_ready;
  wire [27:0] extsi92_outs;
  wire  extsi92_outs_valid;
  wire  extsi92_outs_ready;
  wire [24:0] extsi93_outs;
  wire  extsi93_outs_valid;
  wire  extsi93_outs_ready;
  wire [21:0] extsi94_outs;
  wire  extsi94_outs_valid;
  wire  extsi94_outs_ready;
  wire [18:0] extsi95_outs;
  wire  extsi95_outs_valid;
  wire  extsi95_outs_ready;
  wire [15:0] extsi96_outs;
  wire  extsi96_outs_valid;
  wire  extsi96_outs_ready;
  wire [11:0] extsi97_outs;
  wire  extsi97_outs_valid;
  wire  extsi97_outs_ready;
  wire  source19_outs_valid;
  wire  source19_outs_ready;
  wire [3:0] constant261_outs;
  wire  constant261_outs_valid;
  wire  constant261_outs_ready;
  wire [12:0] extui0_outs;
  wire  extui0_outs_valid;
  wire  extui0_outs_ready;
  wire [12:0] extsi145_outs;
  wire  extsi145_outs_valid;
  wire  extsi145_outs_ready;
  wire [15:0] extsi146_outs;
  wire  extsi146_outs_valid;
  wire  extsi146_outs_ready;
  wire [19:0] extsi147_outs;
  wire  extsi147_outs_valid;
  wire  extsi147_outs_ready;
  wire [22:0] extsi148_outs;
  wire  extsi148_outs_valid;
  wire  extsi148_outs_ready;
  wire [25:0] extsi149_outs;
  wire  extsi149_outs_valid;
  wire  extsi149_outs_ready;
  wire [28:0] extsi150_outs;
  wire  extsi150_outs_valid;
  wire  extsi150_outs_ready;
  wire [31:0] extsi151_outs;
  wire  extsi151_outs_valid;
  wire  extsi151_outs_ready;
  wire [34:0] extsi152_outs;
  wire  extsi152_outs_valid;
  wire  extsi152_outs_ready;
  wire [37:0] extsi153_outs;
  wire  extsi153_outs_valid;
  wire  extsi153_outs_ready;
  wire [41:0] extsi154_outs;
  wire  extsi154_outs_valid;
  wire  extsi154_outs_ready;
  wire [12:0] muli0_result;
  wire  muli0_result_valid;
  wire  muli0_result_ready;
  wire [10:0] trunci2_outs;
  wire  trunci2_outs_valid;
  wire  trunci2_outs_ready;
  wire [7:0] buffer60_outs;
  wire  buffer60_outs_valid;
  wire  buffer60_outs_ready;
  wire [7:0] buffer61_outs;
  wire  buffer61_outs_valid;
  wire  buffer61_outs_ready;
  wire [11:0] extsi3_outs;
  wire  extsi3_outs_valid;
  wire  extsi3_outs_ready;
  wire [11:0] shli0_result;
  wire  shli0_result_valid;
  wire  shli0_result_ready;
  wire [10:0] trunci24_outs;
  wire  trunci24_outs_valid;
  wire  trunci24_outs_ready;
  wire [10:0] addi0_result;
  wire  addi0_result_valid;
  wire  addi0_result_ready;
  wire [15:0] extsi155_outs;
  wire  extsi155_outs_valid;
  wire  extsi155_outs_ready;
  wire [15:0] muli1_result;
  wire  muli1_result_valid;
  wire  muli1_result_ready;
  wire [14:0] trunci4_outs;
  wire  trunci4_outs_valid;
  wire  trunci4_outs_ready;
  wire [11:0] buffer58_outs;
  wire  buffer58_outs_valid;
  wire  buffer58_outs_ready;
  wire [11:0] buffer59_outs;
  wire  buffer59_outs_valid;
  wire  buffer59_outs_ready;
  wire [15:0] extsi7_outs;
  wire  extsi7_outs_valid;
  wire  extsi7_outs_ready;
  wire [15:0] shli1_result;
  wire  shli1_result_valid;
  wire  shli1_result_ready;
  wire [14:0] trunci25_outs;
  wire  trunci25_outs_valid;
  wire  trunci25_outs_ready;
  wire [14:0] addi1_result;
  wire  addi1_result_valid;
  wire  addi1_result_ready;
  wire [19:0] extsi156_outs;
  wire  extsi156_outs_valid;
  wire  extsi156_outs_ready;
  wire [19:0] muli2_result;
  wire  muli2_result_valid;
  wire  muli2_result_ready;
  wire [17:0] trunci6_outs;
  wire  trunci6_outs_valid;
  wire  trunci6_outs_ready;
  wire [13:0] buffer56_outs;
  wire  buffer56_outs_valid;
  wire  buffer56_outs_ready;
  wire [13:0] buffer57_outs;
  wire  buffer57_outs_valid;
  wire  buffer57_outs_ready;
  wire [18:0] extsi11_outs;
  wire  extsi11_outs_valid;
  wire  extsi11_outs_ready;
  wire [18:0] shli2_result;
  wire  shli2_result_valid;
  wire  shli2_result_ready;
  wire [17:0] trunci26_outs;
  wire  trunci26_outs_valid;
  wire  trunci26_outs_ready;
  wire [17:0] addi2_result;
  wire  addi2_result_valid;
  wire  addi2_result_ready;
  wire [22:0] extsi157_outs;
  wire  extsi157_outs_valid;
  wire  extsi157_outs_ready;
  wire [22:0] muli3_result;
  wire  muli3_result_valid;
  wire  muli3_result_ready;
  wire [20:0] trunci8_outs;
  wire  trunci8_outs_valid;
  wire  trunci8_outs_ready;
  wire [17:0] buffer54_outs;
  wire  buffer54_outs_valid;
  wire  buffer54_outs_ready;
  wire [17:0] buffer55_outs;
  wire  buffer55_outs_valid;
  wire  buffer55_outs_ready;
  wire [21:0] extsi15_outs;
  wire  extsi15_outs_valid;
  wire  extsi15_outs_ready;
  wire [21:0] shli3_result;
  wire  shli3_result_valid;
  wire  shli3_result_ready;
  wire [20:0] trunci27_outs;
  wire  trunci27_outs_valid;
  wire  trunci27_outs_ready;
  wire [20:0] addi3_result;
  wire  addi3_result_valid;
  wire  addi3_result_ready;
  wire [25:0] extsi158_outs;
  wire  extsi158_outs_valid;
  wire  extsi158_outs_ready;
  wire [25:0] muli4_result;
  wire  muli4_result_valid;
  wire  muli4_result_ready;
  wire [23:0] trunci10_outs;
  wire  trunci10_outs_valid;
  wire  trunci10_outs_ready;
  wire [20:0] buffer52_outs;
  wire  buffer52_outs_valid;
  wire  buffer52_outs_ready;
  wire [20:0] buffer53_outs;
  wire  buffer53_outs_valid;
  wire  buffer53_outs_ready;
  wire [24:0] extsi19_outs;
  wire  extsi19_outs_valid;
  wire  extsi19_outs_ready;
  wire [24:0] shli4_result;
  wire  shli4_result_valid;
  wire  shli4_result_ready;
  wire [23:0] trunci28_outs;
  wire  trunci28_outs_valid;
  wire  trunci28_outs_ready;
  wire [23:0] addi4_result;
  wire  addi4_result_valid;
  wire  addi4_result_ready;
  wire [28:0] extsi159_outs;
  wire  extsi159_outs_valid;
  wire  extsi159_outs_ready;
  wire [28:0] muli5_result;
  wire  muli5_result_valid;
  wire  muli5_result_ready;
  wire [26:0] trunci12_outs;
  wire  trunci12_outs_valid;
  wire  trunci12_outs_ready;
  wire [23:0] buffer50_outs;
  wire  buffer50_outs_valid;
  wire  buffer50_outs_ready;
  wire [23:0] buffer51_outs;
  wire  buffer51_outs_valid;
  wire  buffer51_outs_ready;
  wire [27:0] extsi23_outs;
  wire  extsi23_outs_valid;
  wire  extsi23_outs_ready;
  wire [27:0] shli5_result;
  wire  shli5_result_valid;
  wire  shli5_result_ready;
  wire [26:0] trunci29_outs;
  wire  trunci29_outs_valid;
  wire  trunci29_outs_ready;
  wire [26:0] addi5_result;
  wire  addi5_result_valid;
  wire  addi5_result_ready;
  wire [31:0] extsi160_outs;
  wire  extsi160_outs_valid;
  wire  extsi160_outs_ready;
  wire [31:0] muli6_result;
  wire  muli6_result_valid;
  wire  muli6_result_ready;
  wire [29:0] trunci14_outs;
  wire  trunci14_outs_valid;
  wire  trunci14_outs_ready;
  wire [26:0] buffer48_outs;
  wire  buffer48_outs_valid;
  wire  buffer48_outs_ready;
  wire [26:0] buffer49_outs;
  wire  buffer49_outs_valid;
  wire  buffer49_outs_ready;
  wire [30:0] extsi27_outs;
  wire  extsi27_outs_valid;
  wire  extsi27_outs_ready;
  wire [30:0] shli6_result;
  wire  shli6_result_valid;
  wire  shli6_result_ready;
  wire [29:0] trunci30_outs;
  wire  trunci30_outs_valid;
  wire  trunci30_outs_ready;
  wire [29:0] addi6_result;
  wire  addi6_result_valid;
  wire  addi6_result_ready;
  wire [34:0] extsi161_outs;
  wire  extsi161_outs_valid;
  wire  extsi161_outs_ready;
  wire [34:0] muli7_result;
  wire  muli7_result_valid;
  wire  muli7_result_ready;
  wire [32:0] trunci16_outs;
  wire  trunci16_outs_valid;
  wire  trunci16_outs_ready;
  wire [29:0] buffer46_outs;
  wire  buffer46_outs_valid;
  wire  buffer46_outs_ready;
  wire [29:0] buffer47_outs;
  wire  buffer47_outs_valid;
  wire  buffer47_outs_ready;
  wire [33:0] extsi31_outs;
  wire  extsi31_outs_valid;
  wire  extsi31_outs_ready;
  wire [33:0] shli7_result;
  wire  shli7_result_valid;
  wire  shli7_result_ready;
  wire [32:0] trunci31_outs;
  wire  trunci31_outs_valid;
  wire  trunci31_outs_ready;
  wire [32:0] addi7_result;
  wire  addi7_result_valid;
  wire  addi7_result_ready;
  wire [37:0] extsi162_outs;
  wire  extsi162_outs_valid;
  wire  extsi162_outs_ready;
  wire [37:0] muli8_result;
  wire  muli8_result_valid;
  wire  muli8_result_ready;
  wire [36:0] trunci18_outs;
  wire  trunci18_outs_valid;
  wire  trunci18_outs_ready;
  wire [33:0] buffer44_outs;
  wire  buffer44_outs_valid;
  wire  buffer44_outs_ready;
  wire [33:0] buffer45_outs;
  wire  buffer45_outs_valid;
  wire  buffer45_outs_ready;
  wire [37:0] extsi35_outs;
  wire  extsi35_outs_valid;
  wire  extsi35_outs_ready;
  wire [37:0] shli8_result;
  wire  shli8_result_valid;
  wire  shli8_result_ready;
  wire [36:0] trunci32_outs;
  wire  trunci32_outs_valid;
  wire  trunci32_outs_ready;
  wire [36:0] addi8_result;
  wire  addi8_result_valid;
  wire  addi8_result_ready;
  wire [41:0] extsi163_outs;
  wire  extsi163_outs_valid;
  wire  extsi163_outs_ready;
  wire [41:0] muli9_result;
  wire  muli9_result_valid;
  wire  muli9_result_ready;
  wire [12:0] trunci33_outs;
  wire  trunci33_outs_valid;
  wire  trunci33_outs_ready;
  wire [35:0] buffer42_outs;
  wire  buffer42_outs_valid;
  wire  buffer42_outs_ready;
  wire [35:0] buffer43_outs;
  wire  buffer43_outs_valid;
  wire  buffer43_outs_ready;
  wire [39:0] extsi39_outs;
  wire  extsi39_outs_valid;
  wire  extsi39_outs_ready;
  wire [39:0] shli9_result;
  wire  shli9_result_valid;
  wire  shli9_result_ready;
  wire [12:0] trunci34_outs;
  wire  trunci34_outs_valid;
  wire  trunci34_outs_ready;
  wire [12:0] addi9_result;
  wire  addi9_result_valid;
  wire  addi9_result_ready;
  wire [12:0] shrsi0_result;
  wire  shrsi0_result_valid;
  wire  shrsi0_result_ready;
  wire [7:0] trunci22_outs;
  wire  trunci22_outs_valid;
  wire  trunci22_outs_ready;

  assign out0 = trunci22_outs;
  assign out0_valid = trunci22_outs_valid;
  assign trunci22_outs_ready = out0_ready;
  assign end_valid = fork0_outs_11_valid;
  assign fork0_outs_11_ready = end_ready;

  fork_dataless #(.SIZE(13)) fork0(
    .ins_valid (start_valid),
    .ins_ready (start_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork0_outs_12_valid, fork0_outs_11_valid, fork0_outs_10_valid, fork0_outs_9_valid, fork0_outs_8_valid, fork0_outs_7_valid, fork0_outs_6_valid, fork0_outs_5_valid, fork0_outs_4_valid, fork0_outs_3_valid, fork0_outs_2_valid, fork0_outs_1_valid, fork0_outs_0_valid}),
    .outs_ready ({fork0_outs_12_ready, fork0_outs_11_ready, fork0_outs_10_ready, fork0_outs_9_ready, fork0_outs_8_ready, fork0_outs_7_ready, fork0_outs_6_ready, fork0_outs_5_ready, fork0_outs_4_ready, fork0_outs_3_ready, fork0_outs_2_ready, fork0_outs_1_ready, fork0_outs_0_ready})
  );

  fork_type #(.SIZE(2), .DATA_TYPE(8)) fork1(
    .ins (in0),
    .ins_valid (in0_valid),
    .ins_ready (in0_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork1_outs_1, fork1_outs_0}),
    .outs_valid ({fork1_outs_1_valid, fork1_outs_0_valid}),
    .outs_ready ({fork1_outs_1_ready, fork1_outs_0_ready})
  );

  trunci #(.INPUT_TYPE(8), .OUTPUT_TYPE(5)) trunci23(
    .ins (fork1_outs_0),
    .ins_valid (fork1_outs_0_valid),
    .ins_ready (fork1_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci23_outs),
    .outs_valid (trunci23_outs_valid),
    .outs_ready (trunci23_outs_ready)
  );

  source source0(
    .clk (clk),
    .rst (rst),
    .outs_valid (source0_outs_valid),
    .outs_ready (source0_outs_ready)
  );

  handshake_constant_0 #(.DATA_WIDTH(1)) constant212(
    .ctrl_valid (source0_outs_valid),
    .ctrl_ready (source0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant212_outs),
    .outs_valid (constant212_outs_valid),
    .outs_ready (constant212_outs_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(3)) extsi99(
    .ins (constant212_outs),
    .ins_valid (constant212_outs_valid),
    .ins_ready (constant212_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi99_outs),
    .outs_valid (extsi99_outs_valid),
    .outs_ready (extsi99_outs_ready)
  );

  handshake_constant_1 #(.DATA_WIDTH(8)) constant94(
    .ctrl_valid (fork0_outs_10_valid),
    .ctrl_ready (fork0_outs_10_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant94_outs),
    .outs_valid (constant94_outs_valid),
    .outs_ready (constant94_outs_ready)
  );

  handshake_constant_2 #(.DATA_WIDTH(7)) constant213(
    .ctrl_valid (fork0_outs_1_valid),
    .ctrl_ready (fork0_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant213_outs),
    .outs_valid (constant213_outs_valid),
    .outs_ready (constant213_outs_ready)
  );

  handshake_constant_3 #(.DATA_WIDTH(12)) constant96(
    .ctrl_valid (fork0_outs_9_valid),
    .ctrl_ready (fork0_outs_9_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant96_outs),
    .outs_valid (constant96_outs_valid),
    .outs_ready (constant96_outs_ready)
  );

  handshake_constant_4 #(.DATA_WIDTH(14)) constant97(
    .ctrl_valid (fork0_outs_8_valid),
    .ctrl_ready (fork0_outs_8_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant97_outs),
    .outs_valid (constant97_outs_valid),
    .outs_ready (constant97_outs_ready)
  );

  handshake_constant_5 #(.DATA_WIDTH(18)) constant98(
    .ctrl_valid (fork0_outs_7_valid),
    .ctrl_ready (fork0_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant98_outs),
    .outs_valid (constant98_outs_valid),
    .outs_ready (constant98_outs_ready)
  );

  handshake_constant_6 #(.DATA_WIDTH(21)) constant99(
    .ctrl_valid (fork0_outs_6_valid),
    .ctrl_ready (fork0_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant99_outs),
    .outs_valid (constant99_outs_valid),
    .outs_ready (constant99_outs_ready)
  );

  handshake_constant_7 #(.DATA_WIDTH(24)) constant100(
    .ctrl_valid (fork0_outs_5_valid),
    .ctrl_ready (fork0_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant100_outs),
    .outs_valid (constant100_outs_valid),
    .outs_ready (constant100_outs_ready)
  );

  handshake_constant_8 #(.DATA_WIDTH(27)) constant101(
    .ctrl_valid (fork0_outs_4_valid),
    .ctrl_ready (fork0_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant101_outs),
    .outs_valid (constant101_outs_valid),
    .outs_ready (constant101_outs_ready)
  );

  handshake_constant_9 #(.DATA_WIDTH(30)) constant102(
    .ctrl_valid (fork0_outs_3_valid),
    .ctrl_ready (fork0_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant102_outs),
    .outs_valid (constant102_outs_valid),
    .outs_ready (constant102_outs_ready)
  );

  handshake_constant_10 #(.DATA_WIDTH(34)) constant103(
    .ctrl_valid (fork0_outs_2_valid),
    .ctrl_ready (fork0_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant103_outs),
    .outs_valid (constant103_outs_valid),
    .outs_ready (constant103_outs_ready)
  );

  handshake_constant_11 #(.DATA_WIDTH(34)) constant214(
    .ctrl_valid (fork0_outs_0_valid),
    .ctrl_ready (fork0_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant214_outs),
    .outs_valid (constant214_outs_valid),
    .outs_ready (constant214_outs_ready)
  );

  source source1(
    .clk (clk),
    .rst (rst),
    .outs_valid (source1_outs_valid),
    .outs_ready (source1_outs_ready)
  );

  handshake_constant_12 #(.DATA_WIDTH(4)) constant215(
    .ctrl_valid (source1_outs_valid),
    .ctrl_ready (source1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant215_outs),
    .outs_valid (constant215_outs_valid),
    .outs_ready (constant215_outs_ready)
  );

  extsi #(.INPUT_TYPE(4), .OUTPUT_TYPE(8)) extsi43(
    .ins (constant215_outs),
    .ins_valid (constant215_outs_valid),
    .ins_ready (constant215_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi43_outs),
    .outs_valid (extsi43_outs_valid),
    .outs_ready (extsi43_outs_ready)
  );

  shrui #(.DATA_TYPE(8)) shrui0(
    .lhs (fork1_outs_1),
    .lhs_valid (fork1_outs_1_valid),
    .lhs_ready (fork1_outs_1_ready),
    .rhs (extsi43_outs),
    .rhs_valid (extsi43_outs_valid),
    .rhs_ready (extsi43_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shrui0_result),
    .result_valid (shrui0_result_valid),
    .result_ready (shrui0_result_ready)
  );

  trunci #(.INPUT_TYPE(8), .OUTPUT_TYPE(3)) trunci0(
    .ins (shrui0_result),
    .ins_valid (shrui0_result_valid),
    .ins_ready (shrui0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci0_outs),
    .outs_valid (trunci0_outs_valid),
    .outs_ready (trunci0_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(3)) fork2(
    .ins (trunci0_outs),
    .ins_valid (trunci0_outs_valid),
    .ins_ready (trunci0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork2_outs_1, fork2_outs_0}),
    .outs_valid ({fork2_outs_1_valid, fork2_outs_0_valid}),
    .outs_ready ({fork2_outs_1_ready, fork2_outs_0_ready})
  );

  handshake_cmpi_0 #(.DATA_TYPE(3)) cmpi0(
    .lhs (fork2_outs_0),
    .lhs_valid (fork2_outs_0_valid),
    .lhs_ready (fork2_outs_0_ready),
    .rhs (extsi99_outs),
    .rhs_valid (extsi99_outs_valid),
    .rhs_ready (extsi99_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi0_result),
    .result_valid (cmpi0_result_valid),
    .result_ready (cmpi0_result_ready)
  );

  fork_type #(.SIZE(14), .DATA_TYPE(1)) fork3(
    .ins (cmpi0_result),
    .ins_valid (cmpi0_result_valid),
    .ins_ready (cmpi0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork3_outs_13, fork3_outs_12, fork3_outs_11, fork3_outs_10, fork3_outs_9, fork3_outs_8, fork3_outs_7, fork3_outs_6, fork3_outs_5, fork3_outs_4, fork3_outs_3, fork3_outs_2, fork3_outs_1, fork3_outs_0}),
    .outs_valid ({fork3_outs_13_valid, fork3_outs_12_valid, fork3_outs_11_valid, fork3_outs_10_valid, fork3_outs_9_valid, fork3_outs_8_valid, fork3_outs_7_valid, fork3_outs_6_valid, fork3_outs_5_valid, fork3_outs_4_valid, fork3_outs_3_valid, fork3_outs_2_valid, fork3_outs_1_valid, fork3_outs_0_valid}),
    .outs_ready ({fork3_outs_13_ready, fork3_outs_12_ready, fork3_outs_11_ready, fork3_outs_10_ready, fork3_outs_9_ready, fork3_outs_8_ready, fork3_outs_7_ready, fork3_outs_6_ready, fork3_outs_5_ready, fork3_outs_4_ready, fork3_outs_3_ready, fork3_outs_2_ready, fork3_outs_1_ready, fork3_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(34)) cond_br8(
    .condition (fork3_outs_13),
    .condition_valid (fork3_outs_13_valid),
    .condition_ready (fork3_outs_13_ready),
    .data (constant214_outs),
    .data_valid (constant214_outs_valid),
    .data_ready (constant214_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br8_trueOut),
    .trueOut_valid (cond_br8_trueOut_valid),
    .trueOut_ready (cond_br8_trueOut_ready),
    .falseOut (cond_br8_falseOut),
    .falseOut_valid (cond_br8_falseOut_valid),
    .falseOut_ready (cond_br8_falseOut_ready)
  );

  sink #(.DATA_TYPE(34)) sink0(
    .ins (cond_br8_falseOut),
    .ins_valid (cond_br8_falseOut_valid),
    .ins_ready (cond_br8_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(34), .OUTPUT_TYPE(36)) extsi100(
    .ins (cond_br8_trueOut),
    .ins_valid (cond_br8_trueOut_valid),
    .ins_ready (cond_br8_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi100_outs),
    .outs_valid (extsi100_outs_valid),
    .outs_ready (extsi100_outs_ready)
  );

  cond_br #(.DATA_TYPE(34)) cond_br9(
    .condition (fork3_outs_10),
    .condition_valid (fork3_outs_10_valid),
    .condition_ready (fork3_outs_10_ready),
    .data (constant103_outs),
    .data_valid (constant103_outs_valid),
    .data_ready (constant103_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br9_trueOut),
    .trueOut_valid (cond_br9_trueOut_valid),
    .trueOut_ready (cond_br9_trueOut_ready),
    .falseOut (cond_br9_falseOut),
    .falseOut_valid (cond_br9_falseOut_valid),
    .falseOut_ready (cond_br9_falseOut_ready)
  );

  sink #(.DATA_TYPE(34)) sink1(
    .ins (cond_br9_falseOut),
    .ins_valid (cond_br9_falseOut_valid),
    .ins_ready (cond_br9_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(30)) cond_br10(
    .condition (fork3_outs_9),
    .condition_valid (fork3_outs_9_valid),
    .condition_ready (fork3_outs_9_ready),
    .data (constant102_outs),
    .data_valid (constant102_outs_valid),
    .data_ready (constant102_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br10_trueOut),
    .trueOut_valid (cond_br10_trueOut_valid),
    .trueOut_ready (cond_br10_trueOut_ready),
    .falseOut (cond_br10_falseOut),
    .falseOut_valid (cond_br10_falseOut_valid),
    .falseOut_ready (cond_br10_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink2(
    .ins (cond_br10_falseOut),
    .ins_valid (cond_br10_falseOut_valid),
    .ins_ready (cond_br10_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br11(
    .condition (fork3_outs_8),
    .condition_valid (fork3_outs_8_valid),
    .condition_ready (fork3_outs_8_ready),
    .data (constant101_outs),
    .data_valid (constant101_outs_valid),
    .data_ready (constant101_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br11_trueOut),
    .trueOut_valid (cond_br11_trueOut_valid),
    .trueOut_ready (cond_br11_trueOut_ready),
    .falseOut (cond_br11_falseOut),
    .falseOut_valid (cond_br11_falseOut_valid),
    .falseOut_ready (cond_br11_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink3(
    .ins (cond_br11_falseOut),
    .ins_valid (cond_br11_falseOut_valid),
    .ins_ready (cond_br11_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(24)) cond_br12(
    .condition (fork3_outs_7),
    .condition_valid (fork3_outs_7_valid),
    .condition_ready (fork3_outs_7_ready),
    .data (constant100_outs),
    .data_valid (constant100_outs_valid),
    .data_ready (constant100_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br12_trueOut),
    .trueOut_valid (cond_br12_trueOut_valid),
    .trueOut_ready (cond_br12_trueOut_ready),
    .falseOut (cond_br12_falseOut),
    .falseOut_valid (cond_br12_falseOut_valid),
    .falseOut_ready (cond_br12_falseOut_ready)
  );

  sink #(.DATA_TYPE(24)) sink4(
    .ins (cond_br12_falseOut),
    .ins_valid (cond_br12_falseOut_valid),
    .ins_ready (cond_br12_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(21)) cond_br13(
    .condition (fork3_outs_6),
    .condition_valid (fork3_outs_6_valid),
    .condition_ready (fork3_outs_6_ready),
    .data (constant99_outs),
    .data_valid (constant99_outs_valid),
    .data_ready (constant99_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br13_trueOut),
    .trueOut_valid (cond_br13_trueOut_valid),
    .trueOut_ready (cond_br13_trueOut_ready),
    .falseOut (cond_br13_falseOut),
    .falseOut_valid (cond_br13_falseOut_valid),
    .falseOut_ready (cond_br13_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink5(
    .ins (cond_br13_falseOut),
    .ins_valid (cond_br13_falseOut_valid),
    .ins_ready (cond_br13_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(18)) cond_br14(
    .condition (fork3_outs_5),
    .condition_valid (fork3_outs_5_valid),
    .condition_ready (fork3_outs_5_ready),
    .data (constant98_outs),
    .data_valid (constant98_outs_valid),
    .data_ready (constant98_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br14_trueOut),
    .trueOut_valid (cond_br14_trueOut_valid),
    .trueOut_ready (cond_br14_trueOut_ready),
    .falseOut (cond_br14_falseOut),
    .falseOut_valid (cond_br14_falseOut_valid),
    .falseOut_ready (cond_br14_falseOut_ready)
  );

  sink #(.DATA_TYPE(18)) sink6(
    .ins (cond_br14_falseOut),
    .ins_valid (cond_br14_falseOut_valid),
    .ins_ready (cond_br14_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(14)) cond_br15(
    .condition (fork3_outs_4),
    .condition_valid (fork3_outs_4_valid),
    .condition_ready (fork3_outs_4_ready),
    .data (constant97_outs),
    .data_valid (constant97_outs_valid),
    .data_ready (constant97_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br15_trueOut),
    .trueOut_valid (cond_br15_trueOut_valid),
    .trueOut_ready (cond_br15_trueOut_ready),
    .falseOut (cond_br15_falseOut),
    .falseOut_valid (cond_br15_falseOut_valid),
    .falseOut_ready (cond_br15_falseOut_ready)
  );

  sink #(.DATA_TYPE(14)) sink7(
    .ins (cond_br15_falseOut),
    .ins_valid (cond_br15_falseOut_valid),
    .ins_ready (cond_br15_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br16(
    .condition (fork3_outs_3),
    .condition_valid (fork3_outs_3_valid),
    .condition_ready (fork3_outs_3_ready),
    .data (constant96_outs),
    .data_valid (constant96_outs_valid),
    .data_ready (constant96_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br16_trueOut),
    .trueOut_valid (cond_br16_trueOut_valid),
    .trueOut_ready (cond_br16_trueOut_ready),
    .falseOut (cond_br16_falseOut),
    .falseOut_valid (cond_br16_falseOut_valid),
    .falseOut_ready (cond_br16_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink8(
    .ins (cond_br16_falseOut),
    .ins_valid (cond_br16_falseOut_valid),
    .ins_ready (cond_br16_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br17(
    .condition (fork3_outs_12),
    .condition_valid (fork3_outs_12_valid),
    .condition_ready (fork3_outs_12_ready),
    .data (constant213_outs),
    .data_valid (constant213_outs_valid),
    .data_ready (constant213_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br17_trueOut),
    .trueOut_valid (cond_br17_trueOut_valid),
    .trueOut_ready (cond_br17_trueOut_ready),
    .falseOut (cond_br17_falseOut),
    .falseOut_valid (cond_br17_falseOut_valid),
    .falseOut_ready (cond_br17_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink9(
    .ins (cond_br17_falseOut),
    .ins_valid (cond_br17_falseOut_valid),
    .ins_ready (cond_br17_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(8)) extsi101(
    .ins (cond_br17_trueOut),
    .ins_valid (cond_br17_trueOut_valid),
    .ins_ready (cond_br17_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi101_outs),
    .outs_valid (extsi101_outs_valid),
    .outs_ready (extsi101_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br18(
    .condition (fork3_outs_2),
    .condition_valid (fork3_outs_2_valid),
    .condition_ready (fork3_outs_2_ready),
    .data (constant94_outs),
    .data_valid (constant94_outs_valid),
    .data_ready (constant94_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br18_trueOut),
    .trueOut_valid (cond_br18_trueOut_valid),
    .trueOut_ready (cond_br18_trueOut_ready),
    .falseOut (cond_br18_falseOut),
    .falseOut_valid (cond_br18_falseOut_valid),
    .falseOut_ready (cond_br18_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink10(
    .ins (cond_br18_falseOut),
    .ins_valid (cond_br18_falseOut_valid),
    .ins_ready (cond_br18_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(5)) cond_br19(
    .condition (fork3_outs_0),
    .condition_valid (fork3_outs_0_valid),
    .condition_ready (fork3_outs_0_ready),
    .data (trunci23_outs),
    .data_valid (trunci23_outs_valid),
    .data_ready (trunci23_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br19_trueOut),
    .trueOut_valid (cond_br19_trueOut_valid),
    .trueOut_ready (cond_br19_trueOut_ready),
    .falseOut (cond_br19_falseOut),
    .falseOut_valid (cond_br19_falseOut_valid),
    .falseOut_ready (cond_br19_falseOut_ready)
  );

  cond_br_dataless cond_br20(
    .condition (fork3_outs_1),
    .condition_valid (fork3_outs_1_valid),
    .condition_ready (fork3_outs_1_ready),
    .data_valid (fork0_outs_12_valid),
    .data_ready (fork0_outs_12_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br20_trueOut_valid),
    .trueOut_ready (cond_br20_trueOut_ready),
    .falseOut_valid (cond_br20_falseOut_valid),
    .falseOut_ready (cond_br20_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(3)) cond_br21(
    .condition (fork3_outs_11),
    .condition_valid (fork3_outs_11_valid),
    .condition_ready (fork3_outs_11_ready),
    .data (fork2_outs_1),
    .data_valid (fork2_outs_1_valid),
    .data_ready (fork2_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br21_trueOut),
    .trueOut_valid (cond_br21_trueOut_valid),
    .trueOut_ready (cond_br21_trueOut_ready),
    .falseOut (cond_br21_falseOut),
    .falseOut_valid (cond_br21_falseOut_valid),
    .falseOut_ready (cond_br21_falseOut_ready)
  );

  sink #(.DATA_TYPE(3)) sink11(
    .ins (cond_br21_trueOut),
    .ins_valid (cond_br21_trueOut_valid),
    .ins_ready (cond_br21_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(3)) buffer2(
    .ins (cond_br21_falseOut),
    .ins_valid (cond_br21_falseOut_valid),
    .ins_ready (cond_br21_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer2_outs),
    .outs_valid (buffer2_outs_valid),
    .outs_ready (buffer2_outs_ready)
  );

  tehb #(.DATA_TYPE(3)) buffer3(
    .ins (buffer2_outs),
    .ins_valid (buffer2_outs_valid),
    .ins_ready (buffer2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer3_outs),
    .outs_valid (buffer3_outs_valid),
    .outs_ready (buffer3_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(3)) fork4(
    .ins (buffer3_outs),
    .ins_valid (buffer3_outs_valid),
    .ins_ready (buffer3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork4_outs_1, fork4_outs_0}),
    .outs_valid ({fork4_outs_1_valid, fork4_outs_0_valid}),
    .outs_ready ({fork4_outs_1_ready, fork4_outs_0_ready})
  );

  oehb_dataless buffer4(
    .ins_valid (cond_br20_falseOut_valid),
    .ins_ready (cond_br20_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer4_outs_valid),
    .outs_ready (buffer4_outs_ready)
  );

  tehb_dataless buffer5(
    .ins_valid (buffer4_outs_valid),
    .ins_ready (buffer4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer5_outs_valid),
    .outs_ready (buffer5_outs_ready)
  );

  fork_dataless #(.SIZE(12)) fork5(
    .ins_valid (buffer5_outs_valid),
    .ins_ready (buffer5_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork5_outs_11_valid, fork5_outs_10_valid, fork5_outs_9_valid, fork5_outs_8_valid, fork5_outs_7_valid, fork5_outs_6_valid, fork5_outs_5_valid, fork5_outs_4_valid, fork5_outs_3_valid, fork5_outs_2_valid, fork5_outs_1_valid, fork5_outs_0_valid}),
    .outs_ready ({fork5_outs_11_ready, fork5_outs_10_ready, fork5_outs_9_ready, fork5_outs_8_ready, fork5_outs_7_ready, fork5_outs_6_ready, fork5_outs_5_ready, fork5_outs_4_ready, fork5_outs_3_ready, fork5_outs_2_ready, fork5_outs_1_ready, fork5_outs_0_ready})
  );

  handshake_constant_13 #(.DATA_WIDTH(35)) constant216(
    .ctrl_valid (fork5_outs_2_valid),
    .ctrl_ready (fork5_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant216_outs),
    .outs_valid (constant216_outs_valid),
    .outs_ready (constant216_outs_ready)
  );

  handshake_constant_14 #(.DATA_WIDTH(33)) constant217(
    .ctrl_valid (fork5_outs_1_valid),
    .ctrl_ready (fork5_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant217_outs),
    .outs_valid (constant217_outs_valid),
    .outs_ready (constant217_outs_ready)
  );

  handshake_constant_15 #(.DATA_WIDTH(30)) constant108(
    .ctrl_valid (fork5_outs_10_valid),
    .ctrl_ready (fork5_outs_10_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant108_outs),
    .outs_valid (constant108_outs_valid),
    .outs_ready (constant108_outs_ready)
  );

  handshake_constant_16 #(.DATA_WIDTH(27)) constant109(
    .ctrl_valid (fork5_outs_9_valid),
    .ctrl_ready (fork5_outs_9_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant109_outs),
    .outs_valid (constant109_outs_valid),
    .outs_ready (constant109_outs_ready)
  );

  handshake_constant_17 #(.DATA_WIDTH(24)) constant110(
    .ctrl_valid (fork5_outs_8_valid),
    .ctrl_ready (fork5_outs_8_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant110_outs),
    .outs_valid (constant110_outs_valid),
    .outs_ready (constant110_outs_ready)
  );

  handshake_constant_18 #(.DATA_WIDTH(21)) constant111(
    .ctrl_valid (fork5_outs_7_valid),
    .ctrl_ready (fork5_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant111_outs),
    .outs_valid (constant111_outs_valid),
    .outs_ready (constant111_outs_ready)
  );

  handshake_constant_19 #(.DATA_WIDTH(18)) constant112(
    .ctrl_valid (fork5_outs_6_valid),
    .ctrl_ready (fork5_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant112_outs),
    .outs_valid (constant112_outs_valid),
    .outs_ready (constant112_outs_ready)
  );

  handshake_constant_20 #(.DATA_WIDTH(14)) constant113(
    .ctrl_valid (fork5_outs_5_valid),
    .ctrl_ready (fork5_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant113_outs),
    .outs_valid (constant113_outs_valid),
    .outs_ready (constant113_outs_ready)
  );

  handshake_constant_21 #(.DATA_WIDTH(9)) constant218(
    .ctrl_valid (fork5_outs_0_valid),
    .ctrl_ready (fork5_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant218_outs),
    .outs_valid (constant218_outs_valid),
    .outs_ready (constant218_outs_ready)
  );

  handshake_constant_22 #(.DATA_WIDTH(8)) constant115(
    .ctrl_valid (fork5_outs_4_valid),
    .ctrl_ready (fork5_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant115_outs),
    .outs_valid (constant115_outs_valid),
    .outs_ready (constant115_outs_ready)
  );

  handshake_constant_23 #(.DATA_WIDTH(8)) constant116(
    .ctrl_valid (fork5_outs_3_valid),
    .ctrl_ready (fork5_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant116_outs),
    .outs_valid (constant116_outs_valid),
    .outs_ready (constant116_outs_ready)
  );

  source source2(
    .clk (clk),
    .rst (rst),
    .outs_valid (source2_outs_valid),
    .outs_ready (source2_outs_ready)
  );

  handshake_constant_24 #(.DATA_WIDTH(2)) constant219(
    .ctrl_valid (source2_outs_valid),
    .ctrl_ready (source2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant219_outs),
    .outs_valid (constant219_outs_valid),
    .outs_ready (constant219_outs_ready)
  );

  extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(3)) extsi102(
    .ins (constant219_outs),
    .ins_valid (constant219_outs_valid),
    .ins_ready (constant219_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi102_outs),
    .outs_valid (extsi102_outs_valid),
    .outs_ready (extsi102_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(3)) cmpi1(
    .lhs (fork4_outs_0),
    .lhs_valid (fork4_outs_0_valid),
    .lhs_ready (fork4_outs_0_ready),
    .rhs (extsi102_outs),
    .rhs_valid (extsi102_outs_valid),
    .rhs_ready (extsi102_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi1_result),
    .result_valid (cmpi1_result_valid),
    .result_ready (cmpi1_result_ready)
  );

  fork_type #(.SIZE(14), .DATA_TYPE(1)) fork6(
    .ins (cmpi1_result),
    .ins_valid (cmpi1_result_valid),
    .ins_ready (cmpi1_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork6_outs_13, fork6_outs_12, fork6_outs_11, fork6_outs_10, fork6_outs_9, fork6_outs_8, fork6_outs_7, fork6_outs_6, fork6_outs_5, fork6_outs_4, fork6_outs_3, fork6_outs_2, fork6_outs_1, fork6_outs_0}),
    .outs_valid ({fork6_outs_13_valid, fork6_outs_12_valid, fork6_outs_11_valid, fork6_outs_10_valid, fork6_outs_9_valid, fork6_outs_8_valid, fork6_outs_7_valid, fork6_outs_6_valid, fork6_outs_5_valid, fork6_outs_4_valid, fork6_outs_3_valid, fork6_outs_2_valid, fork6_outs_1_valid, fork6_outs_0_valid}),
    .outs_ready ({fork6_outs_13_ready, fork6_outs_12_ready, fork6_outs_11_ready, fork6_outs_10_ready, fork6_outs_9_ready, fork6_outs_8_ready, fork6_outs_7_ready, fork6_outs_6_ready, fork6_outs_5_ready, fork6_outs_4_ready, fork6_outs_3_ready, fork6_outs_2_ready, fork6_outs_1_ready, fork6_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(35)) cond_br22(
    .condition (fork6_outs_12),
    .condition_valid (fork6_outs_12_valid),
    .condition_ready (fork6_outs_12_ready),
    .data (constant216_outs),
    .data_valid (constant216_outs_valid),
    .data_ready (constant216_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br22_trueOut),
    .trueOut_valid (cond_br22_trueOut_valid),
    .trueOut_ready (cond_br22_trueOut_ready),
    .falseOut (cond_br22_falseOut),
    .falseOut_valid (cond_br22_falseOut_valid),
    .falseOut_ready (cond_br22_falseOut_ready)
  );

  sink #(.DATA_TYPE(35)) sink13(
    .ins (cond_br22_falseOut),
    .ins_valid (cond_br22_falseOut_valid),
    .ins_ready (cond_br22_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(35), .OUTPUT_TYPE(36)) extsi103(
    .ins (cond_br22_trueOut),
    .ins_valid (cond_br22_trueOut_valid),
    .ins_ready (cond_br22_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi103_outs),
    .outs_valid (extsi103_outs_valid),
    .outs_ready (extsi103_outs_ready)
  );

  cond_br #(.DATA_TYPE(33)) cond_br23(
    .condition (fork6_outs_11),
    .condition_valid (fork6_outs_11_valid),
    .condition_ready (fork6_outs_11_ready),
    .data (constant217_outs),
    .data_valid (constant217_outs_valid),
    .data_ready (constant217_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br23_trueOut),
    .trueOut_valid (cond_br23_trueOut_valid),
    .trueOut_ready (cond_br23_trueOut_ready),
    .falseOut (cond_br23_falseOut),
    .falseOut_valid (cond_br23_falseOut_valid),
    .falseOut_ready (cond_br23_falseOut_ready)
  );

  sink #(.DATA_TYPE(33)) sink14(
    .ins (cond_br23_falseOut),
    .ins_valid (cond_br23_falseOut_valid),
    .ins_ready (cond_br23_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(33), .OUTPUT_TYPE(34)) extsi104(
    .ins (cond_br23_trueOut),
    .ins_valid (cond_br23_trueOut_valid),
    .ins_ready (cond_br23_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi104_outs),
    .outs_valid (extsi104_outs_valid),
    .outs_ready (extsi104_outs_ready)
  );

  cond_br #(.DATA_TYPE(30)) cond_br24(
    .condition (fork6_outs_9),
    .condition_valid (fork6_outs_9_valid),
    .condition_ready (fork6_outs_9_ready),
    .data (constant108_outs),
    .data_valid (constant108_outs_valid),
    .data_ready (constant108_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br24_trueOut),
    .trueOut_valid (cond_br24_trueOut_valid),
    .trueOut_ready (cond_br24_trueOut_ready),
    .falseOut (cond_br24_falseOut),
    .falseOut_valid (cond_br24_falseOut_valid),
    .falseOut_ready (cond_br24_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink15(
    .ins (cond_br24_falseOut),
    .ins_valid (cond_br24_falseOut_valid),
    .ins_ready (cond_br24_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br25(
    .condition (fork6_outs_8),
    .condition_valid (fork6_outs_8_valid),
    .condition_ready (fork6_outs_8_ready),
    .data (constant109_outs),
    .data_valid (constant109_outs_valid),
    .data_ready (constant109_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br25_trueOut),
    .trueOut_valid (cond_br25_trueOut_valid),
    .trueOut_ready (cond_br25_trueOut_ready),
    .falseOut (cond_br25_falseOut),
    .falseOut_valid (cond_br25_falseOut_valid),
    .falseOut_ready (cond_br25_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink16(
    .ins (cond_br25_falseOut),
    .ins_valid (cond_br25_falseOut_valid),
    .ins_ready (cond_br25_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(24)) cond_br26(
    .condition (fork6_outs_7),
    .condition_valid (fork6_outs_7_valid),
    .condition_ready (fork6_outs_7_ready),
    .data (constant110_outs),
    .data_valid (constant110_outs_valid),
    .data_ready (constant110_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br26_trueOut),
    .trueOut_valid (cond_br26_trueOut_valid),
    .trueOut_ready (cond_br26_trueOut_ready),
    .falseOut (cond_br26_falseOut),
    .falseOut_valid (cond_br26_falseOut_valid),
    .falseOut_ready (cond_br26_falseOut_ready)
  );

  sink #(.DATA_TYPE(24)) sink17(
    .ins (cond_br26_falseOut),
    .ins_valid (cond_br26_falseOut_valid),
    .ins_ready (cond_br26_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(21)) cond_br27(
    .condition (fork6_outs_6),
    .condition_valid (fork6_outs_6_valid),
    .condition_ready (fork6_outs_6_ready),
    .data (constant111_outs),
    .data_valid (constant111_outs_valid),
    .data_ready (constant111_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br27_trueOut),
    .trueOut_valid (cond_br27_trueOut_valid),
    .trueOut_ready (cond_br27_trueOut_ready),
    .falseOut (cond_br27_falseOut),
    .falseOut_valid (cond_br27_falseOut_valid),
    .falseOut_ready (cond_br27_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink18(
    .ins (cond_br27_falseOut),
    .ins_valid (cond_br27_falseOut_valid),
    .ins_ready (cond_br27_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(18)) cond_br28(
    .condition (fork6_outs_5),
    .condition_valid (fork6_outs_5_valid),
    .condition_ready (fork6_outs_5_ready),
    .data (constant112_outs),
    .data_valid (constant112_outs_valid),
    .data_ready (constant112_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br28_trueOut),
    .trueOut_valid (cond_br28_trueOut_valid),
    .trueOut_ready (cond_br28_trueOut_ready),
    .falseOut (cond_br28_falseOut),
    .falseOut_valid (cond_br28_falseOut_valid),
    .falseOut_ready (cond_br28_falseOut_ready)
  );

  sink #(.DATA_TYPE(18)) sink19(
    .ins (cond_br28_falseOut),
    .ins_valid (cond_br28_falseOut_valid),
    .ins_ready (cond_br28_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(14)) cond_br29(
    .condition (fork6_outs_4),
    .condition_valid (fork6_outs_4_valid),
    .condition_ready (fork6_outs_4_ready),
    .data (constant113_outs),
    .data_valid (constant113_outs_valid),
    .data_ready (constant113_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br29_trueOut),
    .trueOut_valid (cond_br29_trueOut_valid),
    .trueOut_ready (cond_br29_trueOut_ready),
    .falseOut (cond_br29_falseOut),
    .falseOut_valid (cond_br29_falseOut_valid),
    .falseOut_ready (cond_br29_falseOut_ready)
  );

  sink #(.DATA_TYPE(14)) sink20(
    .ins (cond_br29_falseOut),
    .ins_valid (cond_br29_falseOut_valid),
    .ins_ready (cond_br29_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(9)) cond_br30(
    .condition (fork6_outs_10),
    .condition_valid (fork6_outs_10_valid),
    .condition_ready (fork6_outs_10_ready),
    .data (constant218_outs),
    .data_valid (constant218_outs_valid),
    .data_ready (constant218_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br30_trueOut),
    .trueOut_valid (cond_br30_trueOut_valid),
    .trueOut_ready (cond_br30_trueOut_ready),
    .falseOut (cond_br30_falseOut),
    .falseOut_valid (cond_br30_falseOut_valid),
    .falseOut_ready (cond_br30_falseOut_ready)
  );

  sink #(.DATA_TYPE(9)) sink21(
    .ins (cond_br30_falseOut),
    .ins_valid (cond_br30_falseOut_valid),
    .ins_ready (cond_br30_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(9), .OUTPUT_TYPE(12)) extsi105(
    .ins (cond_br30_trueOut),
    .ins_valid (cond_br30_trueOut_valid),
    .ins_ready (cond_br30_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi105_outs),
    .outs_valid (extsi105_outs_valid),
    .outs_ready (extsi105_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br31(
    .condition (fork6_outs_3),
    .condition_valid (fork6_outs_3_valid),
    .condition_ready (fork6_outs_3_ready),
    .data (constant115_outs),
    .data_valid (constant115_outs_valid),
    .data_ready (constant115_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br31_trueOut),
    .trueOut_valid (cond_br31_trueOut_valid),
    .trueOut_ready (cond_br31_trueOut_ready),
    .falseOut (cond_br31_falseOut),
    .falseOut_valid (cond_br31_falseOut_valid),
    .falseOut_ready (cond_br31_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink22(
    .ins (cond_br31_falseOut),
    .ins_valid (cond_br31_falseOut_valid),
    .ins_ready (cond_br31_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(8)) cond_br32(
    .condition (fork6_outs_2),
    .condition_valid (fork6_outs_2_valid),
    .condition_ready (fork6_outs_2_ready),
    .data (constant116_outs),
    .data_valid (constant116_outs_valid),
    .data_ready (constant116_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br32_trueOut),
    .trueOut_valid (cond_br32_trueOut_valid),
    .trueOut_ready (cond_br32_trueOut_ready),
    .falseOut (cond_br32_falseOut),
    .falseOut_valid (cond_br32_falseOut_valid),
    .falseOut_ready (cond_br32_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink23(
    .ins (cond_br32_falseOut),
    .ins_valid (cond_br32_falseOut_valid),
    .ins_ready (cond_br32_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer0(
    .ins (cond_br19_falseOut),
    .ins_valid (cond_br19_falseOut_valid),
    .ins_ready (cond_br19_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer0_outs),
    .outs_valid (buffer0_outs_valid),
    .outs_ready (buffer0_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer1(
    .ins (buffer0_outs),
    .ins_valid (buffer0_outs_valid),
    .ins_ready (buffer0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer1_outs),
    .outs_valid (buffer1_outs_valid),
    .outs_ready (buffer1_outs_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br33(
    .condition (fork6_outs_0),
    .condition_valid (fork6_outs_0_valid),
    .condition_ready (fork6_outs_0_ready),
    .data (buffer1_outs),
    .data_valid (buffer1_outs_valid),
    .data_ready (buffer1_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br33_trueOut),
    .trueOut_valid (cond_br33_trueOut_valid),
    .trueOut_ready (cond_br33_trueOut_ready),
    .falseOut (cond_br33_falseOut),
    .falseOut_valid (cond_br33_falseOut_valid),
    .falseOut_ready (cond_br33_falseOut_ready)
  );

  cond_br_dataless cond_br34(
    .condition (fork6_outs_1),
    .condition_valid (fork6_outs_1_valid),
    .condition_ready (fork6_outs_1_ready),
    .data_valid (fork5_outs_11_valid),
    .data_ready (fork5_outs_11_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br34_trueOut_valid),
    .trueOut_ready (cond_br34_trueOut_ready),
    .falseOut_valid (cond_br34_falseOut_valid),
    .falseOut_ready (cond_br34_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(3)) cond_br35(
    .condition (fork6_outs_13),
    .condition_valid (fork6_outs_13_valid),
    .condition_ready (fork6_outs_13_ready),
    .data (fork4_outs_1),
    .data_valid (fork4_outs_1_valid),
    .data_ready (fork4_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br35_trueOut),
    .trueOut_valid (cond_br35_trueOut_valid),
    .trueOut_ready (cond_br35_trueOut_ready),
    .falseOut (cond_br35_falseOut),
    .falseOut_valid (cond_br35_falseOut_valid),
    .falseOut_ready (cond_br35_falseOut_ready)
  );

  sink #(.DATA_TYPE(3)) sink24(
    .ins (cond_br35_trueOut),
    .ins_valid (cond_br35_trueOut_valid),
    .ins_ready (cond_br35_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(3)) buffer8(
    .ins (cond_br35_falseOut),
    .ins_valid (cond_br35_falseOut_valid),
    .ins_ready (cond_br35_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer8_outs),
    .outs_valid (buffer8_outs_valid),
    .outs_ready (buffer8_outs_ready)
  );

  tehb #(.DATA_TYPE(3)) buffer9(
    .ins (buffer8_outs),
    .ins_valid (buffer8_outs_valid),
    .ins_ready (buffer8_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer9_outs),
    .outs_valid (buffer9_outs_valid),
    .outs_ready (buffer9_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(3)) fork7(
    .ins (buffer9_outs),
    .ins_valid (buffer9_outs_valid),
    .ins_ready (buffer9_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork7_outs_1, fork7_outs_0}),
    .outs_valid ({fork7_outs_1_valid, fork7_outs_0_valid}),
    .outs_ready ({fork7_outs_1_ready, fork7_outs_0_ready})
  );

  oehb_dataless buffer10(
    .ins_valid (cond_br34_falseOut_valid),
    .ins_ready (cond_br34_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer10_outs_valid),
    .outs_ready (buffer10_outs_ready)
  );

  tehb_dataless buffer11(
    .ins_valid (buffer10_outs_valid),
    .ins_ready (buffer10_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer11_outs_valid),
    .outs_ready (buffer11_outs_ready)
  );

  fork_dataless #(.SIZE(12)) fork8(
    .ins_valid (buffer11_outs_valid),
    .ins_ready (buffer11_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork8_outs_11_valid, fork8_outs_10_valid, fork8_outs_9_valid, fork8_outs_8_valid, fork8_outs_7_valid, fork8_outs_6_valid, fork8_outs_5_valid, fork8_outs_4_valid, fork8_outs_3_valid, fork8_outs_2_valid, fork8_outs_1_valid, fork8_outs_0_valid}),
    .outs_ready ({fork8_outs_11_ready, fork8_outs_10_ready, fork8_outs_9_ready, fork8_outs_8_ready, fork8_outs_7_ready, fork8_outs_6_ready, fork8_outs_5_ready, fork8_outs_4_ready, fork8_outs_3_ready, fork8_outs_2_ready, fork8_outs_1_ready, fork8_outs_0_ready})
  );

  handshake_constant_25 #(.DATA_WIDTH(36)) constant118(
    .ctrl_valid (fork8_outs_10_valid),
    .ctrl_ready (fork8_outs_10_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant118_outs),
    .outs_valid (constant118_outs_valid),
    .outs_ready (constant118_outs_ready)
  );

  handshake_constant_26 #(.DATA_WIDTH(33)) constant220(
    .ctrl_valid (fork8_outs_6_valid),
    .ctrl_ready (fork8_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant220_outs),
    .outs_valid (constant220_outs_valid),
    .outs_ready (constant220_outs_ready)
  );

  handshake_constant_27 #(.DATA_WIDTH(30)) constant120(
    .ctrl_valid (fork8_outs_9_valid),
    .ctrl_ready (fork8_outs_9_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant120_outs),
    .outs_valid (constant120_outs_valid),
    .outs_ready (constant120_outs_ready)
  );

  handshake_constant_28 #(.DATA_WIDTH(26)) constant221(
    .ctrl_valid (fork8_outs_5_valid),
    .ctrl_ready (fork8_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant221_outs),
    .outs_valid (constant221_outs_valid),
    .outs_ready (constant221_outs_ready)
  );

  handshake_constant_29 #(.DATA_WIDTH(22)) constant222(
    .ctrl_valid (fork8_outs_4_valid),
    .ctrl_ready (fork8_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant222_outs),
    .outs_valid (constant222_outs_valid),
    .outs_ready (constant222_outs_ready)
  );

  handshake_constant_30 #(.DATA_WIDTH(21)) constant123(
    .ctrl_valid (fork8_outs_8_valid),
    .ctrl_ready (fork8_outs_8_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant123_outs),
    .outs_valid (constant123_outs_valid),
    .outs_ready (constant123_outs_ready)
  );

  handshake_constant_31 #(.DATA_WIDTH(16)) constant223(
    .ctrl_valid (fork8_outs_3_valid),
    .ctrl_ready (fork8_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant223_outs),
    .outs_valid (constant223_outs_valid),
    .outs_ready (constant223_outs_ready)
  );

  handshake_constant_32 #(.DATA_WIDTH(12)) constant224(
    .ctrl_valid (fork8_outs_2_valid),
    .ctrl_ready (fork8_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant224_outs),
    .outs_valid (constant224_outs_valid),
    .outs_ready (constant224_outs_ready)
  );

  handshake_constant_33 #(.DATA_WIDTH(12)) constant126(
    .ctrl_valid (fork8_outs_7_valid),
    .ctrl_ready (fork8_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant126_outs),
    .outs_valid (constant126_outs_valid),
    .outs_ready (constant126_outs_ready)
  );

  handshake_constant_34 #(.DATA_WIDTH(3)) constant225(
    .ctrl_valid (fork8_outs_1_valid),
    .ctrl_ready (fork8_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant225_outs),
    .outs_valid (constant225_outs_valid),
    .outs_ready (constant225_outs_ready)
  );

  handshake_constant_35 #(.DATA_WIDTH(7)) constant226(
    .ctrl_valid (fork8_outs_0_valid),
    .ctrl_ready (fork8_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant226_outs),
    .outs_valid (constant226_outs_valid),
    .outs_ready (constant226_outs_ready)
  );

  source source3(
    .clk (clk),
    .rst (rst),
    .outs_valid (source3_outs_valid),
    .outs_ready (source3_outs_ready)
  );

  handshake_constant_34 #(.DATA_WIDTH(3)) constant227(
    .ctrl_valid (source3_outs_valid),
    .ctrl_ready (source3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant227_outs),
    .outs_valid (constant227_outs_valid),
    .outs_ready (constant227_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(3)) cmpi2(
    .lhs (fork7_outs_0),
    .lhs_valid (fork7_outs_0_valid),
    .lhs_ready (fork7_outs_0_ready),
    .rhs (constant227_outs),
    .rhs_valid (constant227_outs_valid),
    .rhs_ready (constant227_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi2_result),
    .result_valid (cmpi2_result_valid),
    .result_ready (cmpi2_result_ready)
  );

  fork_type #(.SIZE(14), .DATA_TYPE(1)) fork9(
    .ins (cmpi2_result),
    .ins_valid (cmpi2_result_valid),
    .ins_ready (cmpi2_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork9_outs_13, fork9_outs_12, fork9_outs_11, fork9_outs_10, fork9_outs_9, fork9_outs_8, fork9_outs_7, fork9_outs_6, fork9_outs_5, fork9_outs_4, fork9_outs_3, fork9_outs_2, fork9_outs_1, fork9_outs_0}),
    .outs_valid ({fork9_outs_13_valid, fork9_outs_12_valid, fork9_outs_11_valid, fork9_outs_10_valid, fork9_outs_9_valid, fork9_outs_8_valid, fork9_outs_7_valid, fork9_outs_6_valid, fork9_outs_5_valid, fork9_outs_4_valid, fork9_outs_3_valid, fork9_outs_2_valid, fork9_outs_1_valid, fork9_outs_0_valid}),
    .outs_ready ({fork9_outs_13_ready, fork9_outs_12_ready, fork9_outs_11_ready, fork9_outs_10_ready, fork9_outs_9_ready, fork9_outs_8_ready, fork9_outs_7_ready, fork9_outs_6_ready, fork9_outs_5_ready, fork9_outs_4_ready, fork9_outs_3_ready, fork9_outs_2_ready, fork9_outs_1_ready, fork9_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(36)) cond_br36(
    .condition (fork9_outs_5),
    .condition_valid (fork9_outs_5_valid),
    .condition_ready (fork9_outs_5_ready),
    .data (constant118_outs),
    .data_valid (constant118_outs_valid),
    .data_ready (constant118_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br36_trueOut),
    .trueOut_valid (cond_br36_trueOut_valid),
    .trueOut_ready (cond_br36_trueOut_ready),
    .falseOut (cond_br36_falseOut),
    .falseOut_valid (cond_br36_falseOut_valid),
    .falseOut_ready (cond_br36_falseOut_ready)
  );

  sink #(.DATA_TYPE(36)) sink26(
    .ins (cond_br36_falseOut),
    .ins_valid (cond_br36_falseOut_valid),
    .ins_ready (cond_br36_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(33)) cond_br37(
    .condition (fork9_outs_12),
    .condition_valid (fork9_outs_12_valid),
    .condition_ready (fork9_outs_12_ready),
    .data (constant220_outs),
    .data_valid (constant220_outs_valid),
    .data_ready (constant220_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br37_trueOut),
    .trueOut_valid (cond_br37_trueOut_valid),
    .trueOut_ready (cond_br37_trueOut_ready),
    .falseOut (cond_br37_falseOut),
    .falseOut_valid (cond_br37_falseOut_valid),
    .falseOut_ready (cond_br37_falseOut_ready)
  );

  sink #(.DATA_TYPE(33)) sink27(
    .ins (cond_br37_falseOut),
    .ins_valid (cond_br37_falseOut_valid),
    .ins_ready (cond_br37_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(33), .OUTPUT_TYPE(34)) extsi106(
    .ins (cond_br37_trueOut),
    .ins_valid (cond_br37_trueOut_valid),
    .ins_ready (cond_br37_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi106_outs),
    .outs_valid (extsi106_outs_valid),
    .outs_ready (extsi106_outs_ready)
  );

  cond_br #(.DATA_TYPE(30)) cond_br38(
    .condition (fork9_outs_4),
    .condition_valid (fork9_outs_4_valid),
    .condition_ready (fork9_outs_4_ready),
    .data (constant120_outs),
    .data_valid (constant120_outs_valid),
    .data_ready (constant120_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br38_trueOut),
    .trueOut_valid (cond_br38_trueOut_valid),
    .trueOut_ready (cond_br38_trueOut_ready),
    .falseOut (cond_br38_falseOut),
    .falseOut_valid (cond_br38_falseOut_valid),
    .falseOut_ready (cond_br38_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink28(
    .ins (cond_br38_falseOut),
    .ins_valid (cond_br38_falseOut_valid),
    .ins_ready (cond_br38_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(26)) cond_br39(
    .condition (fork9_outs_11),
    .condition_valid (fork9_outs_11_valid),
    .condition_ready (fork9_outs_11_ready),
    .data (constant221_outs),
    .data_valid (constant221_outs_valid),
    .data_ready (constant221_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br39_trueOut),
    .trueOut_valid (cond_br39_trueOut_valid),
    .trueOut_ready (cond_br39_trueOut_ready),
    .falseOut (cond_br39_falseOut),
    .falseOut_valid (cond_br39_falseOut_valid),
    .falseOut_ready (cond_br39_falseOut_ready)
  );

  sink #(.DATA_TYPE(26)) sink29(
    .ins (cond_br39_falseOut),
    .ins_valid (cond_br39_falseOut_valid),
    .ins_ready (cond_br39_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(26), .OUTPUT_TYPE(27)) extsi107(
    .ins (cond_br39_trueOut),
    .ins_valid (cond_br39_trueOut_valid),
    .ins_ready (cond_br39_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi107_outs),
    .outs_valid (extsi107_outs_valid),
    .outs_ready (extsi107_outs_ready)
  );

  cond_br #(.DATA_TYPE(22)) cond_br40(
    .condition (fork9_outs_10),
    .condition_valid (fork9_outs_10_valid),
    .condition_ready (fork9_outs_10_ready),
    .data (constant222_outs),
    .data_valid (constant222_outs_valid),
    .data_ready (constant222_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br40_trueOut),
    .trueOut_valid (cond_br40_trueOut_valid),
    .trueOut_ready (cond_br40_trueOut_ready),
    .falseOut (cond_br40_falseOut),
    .falseOut_valid (cond_br40_falseOut_valid),
    .falseOut_ready (cond_br40_falseOut_ready)
  );

  sink #(.DATA_TYPE(22)) sink30(
    .ins (cond_br40_falseOut),
    .ins_valid (cond_br40_falseOut_valid),
    .ins_ready (cond_br40_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(22), .OUTPUT_TYPE(24)) extsi108(
    .ins (cond_br40_trueOut),
    .ins_valid (cond_br40_trueOut_valid),
    .ins_ready (cond_br40_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi108_outs),
    .outs_valid (extsi108_outs_valid),
    .outs_ready (extsi108_outs_ready)
  );

  cond_br #(.DATA_TYPE(21)) cond_br41(
    .condition (fork9_outs_3),
    .condition_valid (fork9_outs_3_valid),
    .condition_ready (fork9_outs_3_ready),
    .data (constant123_outs),
    .data_valid (constant123_outs_valid),
    .data_ready (constant123_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br41_trueOut),
    .trueOut_valid (cond_br41_trueOut_valid),
    .trueOut_ready (cond_br41_trueOut_ready),
    .falseOut (cond_br41_falseOut),
    .falseOut_valid (cond_br41_falseOut_valid),
    .falseOut_ready (cond_br41_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink31(
    .ins (cond_br41_falseOut),
    .ins_valid (cond_br41_falseOut_valid),
    .ins_ready (cond_br41_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(16)) cond_br42(
    .condition (fork9_outs_9),
    .condition_valid (fork9_outs_9_valid),
    .condition_ready (fork9_outs_9_ready),
    .data (constant223_outs),
    .data_valid (constant223_outs_valid),
    .data_ready (constant223_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br42_trueOut),
    .trueOut_valid (cond_br42_trueOut_valid),
    .trueOut_ready (cond_br42_trueOut_ready),
    .falseOut (cond_br42_falseOut),
    .falseOut_valid (cond_br42_falseOut_valid),
    .falseOut_ready (cond_br42_falseOut_ready)
  );

  sink #(.DATA_TYPE(16)) sink32(
    .ins (cond_br42_falseOut),
    .ins_valid (cond_br42_falseOut_valid),
    .ins_ready (cond_br42_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(16), .OUTPUT_TYPE(18)) extsi109(
    .ins (cond_br42_trueOut),
    .ins_valid (cond_br42_trueOut_valid),
    .ins_ready (cond_br42_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi109_outs),
    .outs_valid (extsi109_outs_valid),
    .outs_ready (extsi109_outs_ready)
  );

  cond_br #(.DATA_TYPE(12)) cond_br43(
    .condition (fork9_outs_8),
    .condition_valid (fork9_outs_8_valid),
    .condition_ready (fork9_outs_8_ready),
    .data (constant224_outs),
    .data_valid (constant224_outs_valid),
    .data_ready (constant224_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br43_trueOut),
    .trueOut_valid (cond_br43_trueOut_valid),
    .trueOut_ready (cond_br43_trueOut_ready),
    .falseOut (cond_br43_falseOut),
    .falseOut_valid (cond_br43_falseOut_valid),
    .falseOut_ready (cond_br43_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink33(
    .ins (cond_br43_falseOut),
    .ins_valid (cond_br43_falseOut_valid),
    .ins_ready (cond_br43_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(12), .OUTPUT_TYPE(14)) extsi110(
    .ins (cond_br43_trueOut),
    .ins_valid (cond_br43_trueOut_valid),
    .ins_ready (cond_br43_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi110_outs),
    .outs_valid (extsi110_outs_valid),
    .outs_ready (extsi110_outs_ready)
  );

  cond_br #(.DATA_TYPE(12)) cond_br44(
    .condition (fork9_outs_2),
    .condition_valid (fork9_outs_2_valid),
    .condition_ready (fork9_outs_2_ready),
    .data (constant126_outs),
    .data_valid (constant126_outs_valid),
    .data_ready (constant126_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br44_trueOut),
    .trueOut_valid (cond_br44_trueOut_valid),
    .trueOut_ready (cond_br44_trueOut_ready),
    .falseOut (cond_br44_falseOut),
    .falseOut_valid (cond_br44_falseOut_valid),
    .falseOut_ready (cond_br44_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink34(
    .ins (cond_br44_falseOut),
    .ins_valid (cond_br44_falseOut_valid),
    .ins_ready (cond_br44_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(3)) cond_br45(
    .condition (fork9_outs_7),
    .condition_valid (fork9_outs_7_valid),
    .condition_ready (fork9_outs_7_ready),
    .data (constant225_outs),
    .data_valid (constant225_outs_valid),
    .data_ready (constant225_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br45_trueOut),
    .trueOut_valid (cond_br45_trueOut_valid),
    .trueOut_ready (cond_br45_trueOut_ready),
    .falseOut (cond_br45_falseOut),
    .falseOut_valid (cond_br45_falseOut_valid),
    .falseOut_ready (cond_br45_falseOut_ready)
  );

  sink #(.DATA_TYPE(3)) sink35(
    .ins (cond_br45_falseOut),
    .ins_valid (cond_br45_falseOut_valid),
    .ins_ready (cond_br45_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(8)) extsi111(
    .ins (cond_br45_trueOut),
    .ins_valid (cond_br45_trueOut_valid),
    .ins_ready (cond_br45_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi111_outs),
    .outs_valid (extsi111_outs_valid),
    .outs_ready (extsi111_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br46(
    .condition (fork9_outs_6),
    .condition_valid (fork9_outs_6_valid),
    .condition_ready (fork9_outs_6_ready),
    .data (constant226_outs),
    .data_valid (constant226_outs_valid),
    .data_ready (constant226_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br46_trueOut),
    .trueOut_valid (cond_br46_trueOut_valid),
    .trueOut_ready (cond_br46_trueOut_ready),
    .falseOut (cond_br46_falseOut),
    .falseOut_valid (cond_br46_falseOut_valid),
    .falseOut_ready (cond_br46_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink36(
    .ins (cond_br46_falseOut),
    .ins_valid (cond_br46_falseOut_valid),
    .ins_ready (cond_br46_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(8)) extsi112(
    .ins (cond_br46_trueOut),
    .ins_valid (cond_br46_trueOut_valid),
    .ins_ready (cond_br46_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi112_outs),
    .outs_valid (extsi112_outs_valid),
    .outs_ready (extsi112_outs_ready)
  );

  oehb #(.DATA_TYPE(5)) buffer6(
    .ins (cond_br33_falseOut),
    .ins_valid (cond_br33_falseOut_valid),
    .ins_ready (cond_br33_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer6_outs),
    .outs_valid (buffer6_outs_valid),
    .outs_ready (buffer6_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer7(
    .ins (buffer6_outs),
    .ins_valid (buffer6_outs_valid),
    .ins_ready (buffer6_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer7_outs),
    .outs_valid (buffer7_outs_valid),
    .outs_ready (buffer7_outs_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br47(
    .condition (fork9_outs_0),
    .condition_valid (fork9_outs_0_valid),
    .condition_ready (fork9_outs_0_ready),
    .data (buffer7_outs),
    .data_valid (buffer7_outs_valid),
    .data_ready (buffer7_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br47_trueOut),
    .trueOut_valid (cond_br47_trueOut_valid),
    .trueOut_ready (cond_br47_trueOut_ready),
    .falseOut (cond_br47_falseOut),
    .falseOut_valid (cond_br47_falseOut_valid),
    .falseOut_ready (cond_br47_falseOut_ready)
  );

  cond_br_dataless cond_br48(
    .condition (fork9_outs_1),
    .condition_valid (fork9_outs_1_valid),
    .condition_ready (fork9_outs_1_ready),
    .data_valid (fork8_outs_11_valid),
    .data_ready (fork8_outs_11_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br48_trueOut_valid),
    .trueOut_ready (cond_br48_trueOut_ready),
    .falseOut_valid (cond_br48_falseOut_valid),
    .falseOut_ready (cond_br48_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(3)) cond_br49(
    .condition (fork9_outs_13),
    .condition_valid (fork9_outs_13_valid),
    .condition_ready (fork9_outs_13_ready),
    .data (fork7_outs_1),
    .data_valid (fork7_outs_1_valid),
    .data_ready (fork7_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br49_trueOut),
    .trueOut_valid (cond_br49_trueOut_valid),
    .trueOut_ready (cond_br49_trueOut_ready),
    .falseOut (cond_br49_falseOut),
    .falseOut_valid (cond_br49_falseOut_valid),
    .falseOut_ready (cond_br49_falseOut_ready)
  );

  sink #(.DATA_TYPE(3)) sink37(
    .ins (cond_br49_trueOut),
    .ins_valid (cond_br49_trueOut_valid),
    .ins_ready (cond_br49_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(3)) buffer14(
    .ins (cond_br49_falseOut),
    .ins_valid (cond_br49_falseOut_valid),
    .ins_ready (cond_br49_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer14_outs),
    .outs_valid (buffer14_outs_valid),
    .outs_ready (buffer14_outs_ready)
  );

  tehb #(.DATA_TYPE(3)) buffer15(
    .ins (buffer14_outs),
    .ins_valid (buffer14_outs_valid),
    .ins_ready (buffer14_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer15_outs),
    .outs_valid (buffer15_outs_valid),
    .outs_ready (buffer15_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(3)) fork10(
    .ins (buffer15_outs),
    .ins_valid (buffer15_outs_valid),
    .ins_ready (buffer15_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork10_outs_1, fork10_outs_0}),
    .outs_valid ({fork10_outs_1_valid, fork10_outs_0_valid}),
    .outs_ready ({fork10_outs_1_ready, fork10_outs_0_ready})
  );

  oehb_dataless buffer16(
    .ins_valid (cond_br48_falseOut_valid),
    .ins_ready (cond_br48_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer16_outs_valid),
    .outs_ready (buffer16_outs_ready)
  );

  tehb_dataless buffer17(
    .ins_valid (buffer16_outs_valid),
    .ins_ready (buffer16_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer17_outs_valid),
    .outs_ready (buffer17_outs_ready)
  );

  fork_dataless #(.SIZE(12)) fork11(
    .ins_valid (buffer17_outs_valid),
    .ins_ready (buffer17_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork11_outs_11_valid, fork11_outs_10_valid, fork11_outs_9_valid, fork11_outs_8_valid, fork11_outs_7_valid, fork11_outs_6_valid, fork11_outs_5_valid, fork11_outs_4_valid, fork11_outs_3_valid, fork11_outs_2_valid, fork11_outs_1_valid, fork11_outs_0_valid}),
    .outs_ready ({fork11_outs_11_ready, fork11_outs_10_ready, fork11_outs_9_ready, fork11_outs_8_ready, fork11_outs_7_ready, fork11_outs_6_ready, fork11_outs_5_ready, fork11_outs_4_ready, fork11_outs_3_ready, fork11_outs_2_ready, fork11_outs_1_ready, fork11_outs_0_ready})
  );

  handshake_constant_36 #(.DATA_WIDTH(36)) constant130(
    .ctrl_valid (fork11_outs_10_valid),
    .ctrl_ready (fork11_outs_10_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant130_outs),
    .outs_valid (constant130_outs_valid),
    .outs_ready (constant130_outs_ready)
  );

  handshake_constant_37 #(.DATA_WIDTH(32)) constant228(
    .ctrl_valid (fork11_outs_4_valid),
    .ctrl_ready (fork11_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant228_outs),
    .outs_valid (constant228_outs_valid),
    .outs_ready (constant228_outs_ready)
  );

  handshake_constant_38 #(.DATA_WIDTH(30)) constant132(
    .ctrl_valid (fork11_outs_9_valid),
    .ctrl_ready (fork11_outs_9_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant132_outs),
    .outs_valid (constant132_outs_valid),
    .outs_ready (constant132_outs_ready)
  );

  handshake_constant_39 #(.DATA_WIDTH(26)) constant229(
    .ctrl_valid (fork11_outs_3_valid),
    .ctrl_ready (fork11_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant229_outs),
    .outs_valid (constant229_outs_valid),
    .outs_ready (constant229_outs_ready)
  );

  handshake_constant_40 #(.DATA_WIDTH(24)) constant134(
    .ctrl_valid (fork11_outs_8_valid),
    .ctrl_ready (fork11_outs_8_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant134_outs),
    .outs_valid (constant134_outs_valid),
    .outs_ready (constant134_outs_ready)
  );

  handshake_constant_41 #(.DATA_WIDTH(21)) constant135(
    .ctrl_valid (fork11_outs_7_valid),
    .ctrl_ready (fork11_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant135_outs),
    .outs_valid (constant135_outs_valid),
    .outs_ready (constant135_outs_ready)
  );

  handshake_constant_42 #(.DATA_WIDTH(16)) constant230(
    .ctrl_valid (fork11_outs_2_valid),
    .ctrl_ready (fork11_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant230_outs),
    .outs_valid (constant230_outs_valid),
    .outs_ready (constant230_outs_ready)
  );

  handshake_constant_43 #(.DATA_WIDTH(14)) constant137(
    .ctrl_valid (fork11_outs_6_valid),
    .ctrl_ready (fork11_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant137_outs),
    .outs_valid (constant137_outs_valid),
    .outs_ready (constant137_outs_ready)
  );

  handshake_constant_44 #(.DATA_WIDTH(12)) constant138(
    .ctrl_valid (fork11_outs_5_valid),
    .ctrl_ready (fork11_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant138_outs),
    .outs_valid (constant138_outs_valid),
    .outs_ready (constant138_outs_ready)
  );

  handshake_constant_45 #(.DATA_WIDTH(6)) constant231(
    .ctrl_valid (fork11_outs_1_valid),
    .ctrl_ready (fork11_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant231_outs),
    .outs_valid (constant231_outs_valid),
    .outs_ready (constant231_outs_ready)
  );

  handshake_constant_46 #(.DATA_WIDTH(6)) constant232(
    .ctrl_valid (fork11_outs_0_valid),
    .ctrl_ready (fork11_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant232_outs),
    .outs_valid (constant232_outs_valid),
    .outs_ready (constant232_outs_ready)
  );

  source source4(
    .clk (clk),
    .rst (rst),
    .outs_valid (source4_outs_valid),
    .outs_ready (source4_outs_ready)
  );

  handshake_constant_47 #(.DATA_WIDTH(3)) constant233(
    .ctrl_valid (source4_outs_valid),
    .ctrl_ready (source4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant233_outs),
    .outs_valid (constant233_outs_valid),
    .outs_ready (constant233_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(3)) cmpi3(
    .lhs (fork10_outs_0),
    .lhs_valid (fork10_outs_0_valid),
    .lhs_ready (fork10_outs_0_ready),
    .rhs (constant233_outs),
    .rhs_valid (constant233_outs_valid),
    .rhs_ready (constant233_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi3_result),
    .result_valid (cmpi3_result_valid),
    .result_ready (cmpi3_result_ready)
  );

  fork_type #(.SIZE(14), .DATA_TYPE(1)) fork12(
    .ins (cmpi3_result),
    .ins_valid (cmpi3_result_valid),
    .ins_ready (cmpi3_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork12_outs_13, fork12_outs_12, fork12_outs_11, fork12_outs_10, fork12_outs_9, fork12_outs_8, fork12_outs_7, fork12_outs_6, fork12_outs_5, fork12_outs_4, fork12_outs_3, fork12_outs_2, fork12_outs_1, fork12_outs_0}),
    .outs_valid ({fork12_outs_13_valid, fork12_outs_12_valid, fork12_outs_11_valid, fork12_outs_10_valid, fork12_outs_9_valid, fork12_outs_8_valid, fork12_outs_7_valid, fork12_outs_6_valid, fork12_outs_5_valid, fork12_outs_4_valid, fork12_outs_3_valid, fork12_outs_2_valid, fork12_outs_1_valid, fork12_outs_0_valid}),
    .outs_ready ({fork12_outs_13_ready, fork12_outs_12_ready, fork12_outs_11_ready, fork12_outs_10_ready, fork12_outs_9_ready, fork12_outs_8_ready, fork12_outs_7_ready, fork12_outs_6_ready, fork12_outs_5_ready, fork12_outs_4_ready, fork12_outs_3_ready, fork12_outs_2_ready, fork12_outs_1_ready, fork12_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(36)) cond_br50(
    .condition (fork12_outs_7),
    .condition_valid (fork12_outs_7_valid),
    .condition_ready (fork12_outs_7_ready),
    .data (constant130_outs),
    .data_valid (constant130_outs_valid),
    .data_ready (constant130_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br50_trueOut),
    .trueOut_valid (cond_br50_trueOut_valid),
    .trueOut_ready (cond_br50_trueOut_ready),
    .falseOut (cond_br50_falseOut),
    .falseOut_valid (cond_br50_falseOut_valid),
    .falseOut_ready (cond_br50_falseOut_ready)
  );

  sink #(.DATA_TYPE(36)) sink39(
    .ins (cond_br50_falseOut),
    .ins_valid (cond_br50_falseOut_valid),
    .ins_ready (cond_br50_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(32)) cond_br51(
    .condition (fork12_outs_12),
    .condition_valid (fork12_outs_12_valid),
    .condition_ready (fork12_outs_12_ready),
    .data (constant228_outs),
    .data_valid (constant228_outs_valid),
    .data_ready (constant228_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br51_trueOut),
    .trueOut_valid (cond_br51_trueOut_valid),
    .trueOut_ready (cond_br51_trueOut_ready),
    .falseOut (cond_br51_falseOut),
    .falseOut_valid (cond_br51_falseOut_valid),
    .falseOut_ready (cond_br51_falseOut_ready)
  );

  sink #(.DATA_TYPE(32)) sink40(
    .ins (cond_br51_falseOut),
    .ins_valid (cond_br51_falseOut_valid),
    .ins_ready (cond_br51_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(32), .OUTPUT_TYPE(34)) extsi113(
    .ins (cond_br51_trueOut),
    .ins_valid (cond_br51_trueOut_valid),
    .ins_ready (cond_br51_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi113_outs),
    .outs_valid (extsi113_outs_valid),
    .outs_ready (extsi113_outs_ready)
  );

  cond_br #(.DATA_TYPE(30)) cond_br52(
    .condition (fork12_outs_6),
    .condition_valid (fork12_outs_6_valid),
    .condition_ready (fork12_outs_6_ready),
    .data (constant132_outs),
    .data_valid (constant132_outs_valid),
    .data_ready (constant132_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br52_trueOut),
    .trueOut_valid (cond_br52_trueOut_valid),
    .trueOut_ready (cond_br52_trueOut_ready),
    .falseOut (cond_br52_falseOut),
    .falseOut_valid (cond_br52_falseOut_valid),
    .falseOut_ready (cond_br52_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink41(
    .ins (cond_br52_falseOut),
    .ins_valid (cond_br52_falseOut_valid),
    .ins_ready (cond_br52_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(26)) cond_br53(
    .condition (fork12_outs_11),
    .condition_valid (fork12_outs_11_valid),
    .condition_ready (fork12_outs_11_ready),
    .data (constant229_outs),
    .data_valid (constant229_outs_valid),
    .data_ready (constant229_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br53_trueOut),
    .trueOut_valid (cond_br53_trueOut_valid),
    .trueOut_ready (cond_br53_trueOut_ready),
    .falseOut (cond_br53_falseOut),
    .falseOut_valid (cond_br53_falseOut_valid),
    .falseOut_ready (cond_br53_falseOut_ready)
  );

  sink #(.DATA_TYPE(26)) sink42(
    .ins (cond_br53_falseOut),
    .ins_valid (cond_br53_falseOut_valid),
    .ins_ready (cond_br53_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(26), .OUTPUT_TYPE(27)) extsi114(
    .ins (cond_br53_trueOut),
    .ins_valid (cond_br53_trueOut_valid),
    .ins_ready (cond_br53_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi114_outs),
    .outs_valid (extsi114_outs_valid),
    .outs_ready (extsi114_outs_ready)
  );

  cond_br #(.DATA_TYPE(24)) cond_br54(
    .condition (fork12_outs_5),
    .condition_valid (fork12_outs_5_valid),
    .condition_ready (fork12_outs_5_ready),
    .data (constant134_outs),
    .data_valid (constant134_outs_valid),
    .data_ready (constant134_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br54_trueOut),
    .trueOut_valid (cond_br54_trueOut_valid),
    .trueOut_ready (cond_br54_trueOut_ready),
    .falseOut (cond_br54_falseOut),
    .falseOut_valid (cond_br54_falseOut_valid),
    .falseOut_ready (cond_br54_falseOut_ready)
  );

  sink #(.DATA_TYPE(24)) sink43(
    .ins (cond_br54_falseOut),
    .ins_valid (cond_br54_falseOut_valid),
    .ins_ready (cond_br54_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(21)) cond_br55(
    .condition (fork12_outs_4),
    .condition_valid (fork12_outs_4_valid),
    .condition_ready (fork12_outs_4_ready),
    .data (constant135_outs),
    .data_valid (constant135_outs_valid),
    .data_ready (constant135_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br55_trueOut),
    .trueOut_valid (cond_br55_trueOut_valid),
    .trueOut_ready (cond_br55_trueOut_ready),
    .falseOut (cond_br55_falseOut),
    .falseOut_valid (cond_br55_falseOut_valid),
    .falseOut_ready (cond_br55_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink44(
    .ins (cond_br55_falseOut),
    .ins_valid (cond_br55_falseOut_valid),
    .ins_ready (cond_br55_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(16)) cond_br56(
    .condition (fork12_outs_10),
    .condition_valid (fork12_outs_10_valid),
    .condition_ready (fork12_outs_10_ready),
    .data (constant230_outs),
    .data_valid (constant230_outs_valid),
    .data_ready (constant230_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br56_trueOut),
    .trueOut_valid (cond_br56_trueOut_valid),
    .trueOut_ready (cond_br56_trueOut_ready),
    .falseOut (cond_br56_falseOut),
    .falseOut_valid (cond_br56_falseOut_valid),
    .falseOut_ready (cond_br56_falseOut_ready)
  );

  sink #(.DATA_TYPE(16)) sink45(
    .ins (cond_br56_falseOut),
    .ins_valid (cond_br56_falseOut_valid),
    .ins_ready (cond_br56_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(16), .OUTPUT_TYPE(18)) extsi115(
    .ins (cond_br56_trueOut),
    .ins_valid (cond_br56_trueOut_valid),
    .ins_ready (cond_br56_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi115_outs),
    .outs_valid (extsi115_outs_valid),
    .outs_ready (extsi115_outs_ready)
  );

  cond_br #(.DATA_TYPE(14)) cond_br57(
    .condition (fork12_outs_3),
    .condition_valid (fork12_outs_3_valid),
    .condition_ready (fork12_outs_3_ready),
    .data (constant137_outs),
    .data_valid (constant137_outs_valid),
    .data_ready (constant137_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br57_trueOut),
    .trueOut_valid (cond_br57_trueOut_valid),
    .trueOut_ready (cond_br57_trueOut_ready),
    .falseOut (cond_br57_falseOut),
    .falseOut_valid (cond_br57_falseOut_valid),
    .falseOut_ready (cond_br57_falseOut_ready)
  );

  sink #(.DATA_TYPE(14)) sink46(
    .ins (cond_br57_falseOut),
    .ins_valid (cond_br57_falseOut_valid),
    .ins_ready (cond_br57_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br58(
    .condition (fork12_outs_2),
    .condition_valid (fork12_outs_2_valid),
    .condition_ready (fork12_outs_2_ready),
    .data (constant138_outs),
    .data_valid (constant138_outs_valid),
    .data_ready (constant138_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br58_trueOut),
    .trueOut_valid (cond_br58_trueOut_valid),
    .trueOut_ready (cond_br58_trueOut_ready),
    .falseOut (cond_br58_falseOut),
    .falseOut_valid (cond_br58_falseOut_valid),
    .falseOut_ready (cond_br58_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink47(
    .ins (cond_br58_falseOut),
    .ins_valid (cond_br58_falseOut_valid),
    .ins_ready (cond_br58_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(6)) cond_br59(
    .condition (fork12_outs_9),
    .condition_valid (fork12_outs_9_valid),
    .condition_ready (fork12_outs_9_ready),
    .data (constant231_outs),
    .data_valid (constant231_outs_valid),
    .data_ready (constant231_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br59_trueOut),
    .trueOut_valid (cond_br59_trueOut_valid),
    .trueOut_ready (cond_br59_trueOut_ready),
    .falseOut (cond_br59_falseOut),
    .falseOut_valid (cond_br59_falseOut_valid),
    .falseOut_ready (cond_br59_falseOut_ready)
  );

  sink #(.DATA_TYPE(6)) sink48(
    .ins (cond_br59_falseOut),
    .ins_valid (cond_br59_falseOut_valid),
    .ins_ready (cond_br59_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(8)) extsi116(
    .ins (cond_br59_trueOut),
    .ins_valid (cond_br59_trueOut_valid),
    .ins_ready (cond_br59_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi116_outs),
    .outs_valid (extsi116_outs_valid),
    .outs_ready (extsi116_outs_ready)
  );

  cond_br #(.DATA_TYPE(6)) cond_br60(
    .condition (fork12_outs_8),
    .condition_valid (fork12_outs_8_valid),
    .condition_ready (fork12_outs_8_ready),
    .data (constant232_outs),
    .data_valid (constant232_outs_valid),
    .data_ready (constant232_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br60_trueOut),
    .trueOut_valid (cond_br60_trueOut_valid),
    .trueOut_ready (cond_br60_trueOut_ready),
    .falseOut (cond_br60_falseOut),
    .falseOut_valid (cond_br60_falseOut_valid),
    .falseOut_ready (cond_br60_falseOut_ready)
  );

  sink #(.DATA_TYPE(6)) sink49(
    .ins (cond_br60_falseOut),
    .ins_valid (cond_br60_falseOut_valid),
    .ins_ready (cond_br60_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(8)) extsi117(
    .ins (cond_br60_trueOut),
    .ins_valid (cond_br60_trueOut_valid),
    .ins_ready (cond_br60_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi117_outs),
    .outs_valid (extsi117_outs_valid),
    .outs_ready (extsi117_outs_ready)
  );

  oehb #(.DATA_TYPE(5)) buffer12(
    .ins (cond_br47_falseOut),
    .ins_valid (cond_br47_falseOut_valid),
    .ins_ready (cond_br47_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer12_outs),
    .outs_valid (buffer12_outs_valid),
    .outs_ready (buffer12_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer13(
    .ins (buffer12_outs),
    .ins_valid (buffer12_outs_valid),
    .ins_ready (buffer12_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer13_outs),
    .outs_valid (buffer13_outs_valid),
    .outs_ready (buffer13_outs_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br61(
    .condition (fork12_outs_0),
    .condition_valid (fork12_outs_0_valid),
    .condition_ready (fork12_outs_0_ready),
    .data (buffer13_outs),
    .data_valid (buffer13_outs_valid),
    .data_ready (buffer13_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br61_trueOut),
    .trueOut_valid (cond_br61_trueOut_valid),
    .trueOut_ready (cond_br61_trueOut_ready),
    .falseOut (cond_br61_falseOut),
    .falseOut_valid (cond_br61_falseOut_valid),
    .falseOut_ready (cond_br61_falseOut_ready)
  );

  cond_br_dataless cond_br62(
    .condition (fork12_outs_1),
    .condition_valid (fork12_outs_1_valid),
    .condition_ready (fork12_outs_1_ready),
    .data_valid (fork11_outs_11_valid),
    .data_ready (fork11_outs_11_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br62_trueOut_valid),
    .trueOut_ready (cond_br62_trueOut_ready),
    .falseOut_valid (cond_br62_falseOut_valid),
    .falseOut_ready (cond_br62_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(3)) cond_br63(
    .condition (fork12_outs_13),
    .condition_valid (fork12_outs_13_valid),
    .condition_ready (fork12_outs_13_ready),
    .data (fork10_outs_1),
    .data_valid (fork10_outs_1_valid),
    .data_ready (fork10_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br63_trueOut),
    .trueOut_valid (cond_br63_trueOut_valid),
    .trueOut_ready (cond_br63_trueOut_ready),
    .falseOut (cond_br63_falseOut),
    .falseOut_valid (cond_br63_falseOut_valid),
    .falseOut_ready (cond_br63_falseOut_ready)
  );

  sink #(.DATA_TYPE(3)) sink50(
    .ins (cond_br63_trueOut),
    .ins_valid (cond_br63_trueOut_valid),
    .ins_ready (cond_br63_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(3)) buffer20(
    .ins (cond_br63_falseOut),
    .ins_valid (cond_br63_falseOut_valid),
    .ins_ready (cond_br63_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer20_outs),
    .outs_valid (buffer20_outs_valid),
    .outs_ready (buffer20_outs_ready)
  );

  tehb #(.DATA_TYPE(3)) buffer21(
    .ins (buffer20_outs),
    .ins_valid (buffer20_outs_valid),
    .ins_ready (buffer20_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer21_outs),
    .outs_valid (buffer21_outs_valid),
    .outs_ready (buffer21_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(3)) fork13(
    .ins (buffer21_outs),
    .ins_valid (buffer21_outs_valid),
    .ins_ready (buffer21_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork13_outs_1, fork13_outs_0}),
    .outs_valid ({fork13_outs_1_valid, fork13_outs_0_valid}),
    .outs_ready ({fork13_outs_1_ready, fork13_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(4)) extsi118(
    .ins (fork13_outs_0),
    .ins_valid (fork13_outs_0_valid),
    .ins_ready (fork13_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi118_outs),
    .outs_valid (extsi118_outs_valid),
    .outs_ready (extsi118_outs_ready)
  );

  oehb_dataless buffer22(
    .ins_valid (cond_br62_falseOut_valid),
    .ins_ready (cond_br62_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer22_outs_valid),
    .outs_ready (buffer22_outs_ready)
  );

  tehb_dataless buffer23(
    .ins_valid (buffer22_outs_valid),
    .ins_ready (buffer22_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer23_outs_valid),
    .outs_ready (buffer23_outs_ready)
  );

  fork_dataless #(.SIZE(12)) fork14(
    .ins_valid (buffer23_outs_valid),
    .ins_ready (buffer23_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork14_outs_11_valid, fork14_outs_10_valid, fork14_outs_9_valid, fork14_outs_8_valid, fork14_outs_7_valid, fork14_outs_6_valid, fork14_outs_5_valid, fork14_outs_4_valid, fork14_outs_3_valid, fork14_outs_2_valid, fork14_outs_1_valid, fork14_outs_0_valid}),
    .outs_ready ({fork14_outs_11_ready, fork14_outs_10_ready, fork14_outs_9_ready, fork14_outs_8_ready, fork14_outs_7_ready, fork14_outs_6_ready, fork14_outs_5_ready, fork14_outs_4_ready, fork14_outs_3_ready, fork14_outs_2_ready, fork14_outs_1_ready, fork14_outs_0_ready})
  );

  handshake_constant_34 #(.DATA_WIDTH(3)) constant234(
    .ctrl_valid (fork14_outs_5_valid),
    .ctrl_ready (fork14_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant234_outs),
    .outs_valid (constant234_outs_valid),
    .outs_ready (constant234_outs_ready)
  );

  handshake_constant_48 #(.DATA_WIDTH(36)) constant143(
    .ctrl_valid (fork14_outs_10_valid),
    .ctrl_ready (fork14_outs_10_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant143_outs),
    .outs_valid (constant143_outs_valid),
    .outs_ready (constant143_outs_ready)
  );

  handshake_constant_49 #(.DATA_WIDTH(31)) constant235(
    .ctrl_valid (fork14_outs_4_valid),
    .ctrl_ready (fork14_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant235_outs),
    .outs_valid (constant235_outs_valid),
    .outs_ready (constant235_outs_ready)
  );

  handshake_constant_50 #(.DATA_WIDTH(30)) constant145(
    .ctrl_valid (fork14_outs_9_valid),
    .ctrl_ready (fork14_outs_9_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant145_outs),
    .outs_valid (constant145_outs_valid),
    .outs_ready (constant145_outs_ready)
  );

  handshake_constant_51 #(.DATA_WIDTH(25)) constant236(
    .ctrl_valid (fork14_outs_3_valid),
    .ctrl_ready (fork14_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant236_outs),
    .outs_valid (constant236_outs_valid),
    .outs_ready (constant236_outs_ready)
  );

  handshake_constant_52 #(.DATA_WIDTH(24)) constant147(
    .ctrl_valid (fork14_outs_8_valid),
    .ctrl_ready (fork14_outs_8_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant147_outs),
    .outs_valid (constant147_outs_valid),
    .outs_ready (constant147_outs_ready)
  );

  handshake_constant_53 #(.DATA_WIDTH(16)) constant237(
    .ctrl_valid (fork14_outs_2_valid),
    .ctrl_ready (fork14_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant237_outs),
    .outs_valid (constant237_outs_valid),
    .outs_ready (constant237_outs_ready)
  );

  handshake_constant_54 #(.DATA_WIDTH(13)) constant238(
    .ctrl_valid (fork14_outs_1_valid),
    .ctrl_ready (fork14_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant238_outs),
    .outs_valid (constant238_outs_valid),
    .outs_ready (constant238_outs_ready)
  );

  handshake_constant_55 #(.DATA_WIDTH(14)) constant150(
    .ctrl_valid (fork14_outs_7_valid),
    .ctrl_ready (fork14_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant150_outs),
    .outs_valid (constant150_outs_valid),
    .outs_ready (constant150_outs_ready)
  );

  handshake_constant_56 #(.DATA_WIDTH(12)) constant151(
    .ctrl_valid (fork14_outs_6_valid),
    .ctrl_ready (fork14_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant151_outs),
    .outs_valid (constant151_outs_valid),
    .outs_ready (constant151_outs_ready)
  );

  handshake_constant_57 #(.DATA_WIDTH(7)) constant239(
    .ctrl_valid (fork14_outs_0_valid),
    .ctrl_ready (fork14_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant239_outs),
    .outs_valid (constant239_outs_valid),
    .outs_ready (constant239_outs_ready)
  );

  source source5(
    .clk (clk),
    .rst (rst),
    .outs_valid (source5_outs_valid),
    .outs_ready (source5_outs_ready)
  );

  handshake_constant_58 #(.DATA_WIDTH(4)) constant240(
    .ctrl_valid (source5_outs_valid),
    .ctrl_ready (source5_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant240_outs),
    .outs_valid (constant240_outs_valid),
    .outs_ready (constant240_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(4)) cmpi4(
    .lhs (extsi118_outs),
    .lhs_valid (extsi118_outs_valid),
    .lhs_ready (extsi118_outs_ready),
    .rhs (constant240_outs),
    .rhs_valid (constant240_outs_valid),
    .rhs_ready (constant240_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi4_result),
    .result_valid (cmpi4_result_valid),
    .result_ready (cmpi4_result_ready)
  );

  fork_type #(.SIZE(14), .DATA_TYPE(1)) fork15(
    .ins (cmpi4_result),
    .ins_valid (cmpi4_result_valid),
    .ins_ready (cmpi4_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork15_outs_13, fork15_outs_12, fork15_outs_11, fork15_outs_10, fork15_outs_9, fork15_outs_8, fork15_outs_7, fork15_outs_6, fork15_outs_5, fork15_outs_4, fork15_outs_3, fork15_outs_2, fork15_outs_1, fork15_outs_0}),
    .outs_valid ({fork15_outs_13_valid, fork15_outs_12_valid, fork15_outs_11_valid, fork15_outs_10_valid, fork15_outs_9_valid, fork15_outs_8_valid, fork15_outs_7_valid, fork15_outs_6_valid, fork15_outs_5_valid, fork15_outs_4_valid, fork15_outs_3_valid, fork15_outs_2_valid, fork15_outs_1_valid, fork15_outs_0_valid}),
    .outs_ready ({fork15_outs_13_ready, fork15_outs_12_ready, fork15_outs_11_ready, fork15_outs_10_ready, fork15_outs_9_ready, fork15_outs_8_ready, fork15_outs_7_ready, fork15_outs_6_ready, fork15_outs_5_ready, fork15_outs_4_ready, fork15_outs_3_ready, fork15_outs_2_ready, fork15_outs_1_ready, fork15_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(36)) cond_br64(
    .condition (fork15_outs_6),
    .condition_valid (fork15_outs_6_valid),
    .condition_ready (fork15_outs_6_ready),
    .data (constant143_outs),
    .data_valid (constant143_outs_valid),
    .data_ready (constant143_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br64_trueOut),
    .trueOut_valid (cond_br64_trueOut_valid),
    .trueOut_ready (cond_br64_trueOut_ready),
    .falseOut (cond_br64_falseOut),
    .falseOut_valid (cond_br64_falseOut_valid),
    .falseOut_ready (cond_br64_falseOut_ready)
  );

  sink #(.DATA_TYPE(36)) sink52(
    .ins (cond_br64_falseOut),
    .ins_valid (cond_br64_falseOut_valid),
    .ins_ready (cond_br64_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(31)) cond_br65(
    .condition (fork15_outs_12),
    .condition_valid (fork15_outs_12_valid),
    .condition_ready (fork15_outs_12_ready),
    .data (constant235_outs),
    .data_valid (constant235_outs_valid),
    .data_ready (constant235_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br65_trueOut),
    .trueOut_valid (cond_br65_trueOut_valid),
    .trueOut_ready (cond_br65_trueOut_ready),
    .falseOut (cond_br65_falseOut),
    .falseOut_valid (cond_br65_falseOut_valid),
    .falseOut_ready (cond_br65_falseOut_ready)
  );

  sink #(.DATA_TYPE(31)) sink53(
    .ins (cond_br65_falseOut),
    .ins_valid (cond_br65_falseOut_valid),
    .ins_ready (cond_br65_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(31), .OUTPUT_TYPE(34)) extsi119(
    .ins (cond_br65_trueOut),
    .ins_valid (cond_br65_trueOut_valid),
    .ins_ready (cond_br65_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi119_outs),
    .outs_valid (extsi119_outs_valid),
    .outs_ready (extsi119_outs_ready)
  );

  cond_br #(.DATA_TYPE(30)) cond_br66(
    .condition (fork15_outs_5),
    .condition_valid (fork15_outs_5_valid),
    .condition_ready (fork15_outs_5_ready),
    .data (constant145_outs),
    .data_valid (constant145_outs_valid),
    .data_ready (constant145_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br66_trueOut),
    .trueOut_valid (cond_br66_trueOut_valid),
    .trueOut_ready (cond_br66_trueOut_ready),
    .falseOut (cond_br66_falseOut),
    .falseOut_valid (cond_br66_falseOut_valid),
    .falseOut_ready (cond_br66_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink54(
    .ins (cond_br66_falseOut),
    .ins_valid (cond_br66_falseOut_valid),
    .ins_ready (cond_br66_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(25)) cond_br67(
    .condition (fork15_outs_11),
    .condition_valid (fork15_outs_11_valid),
    .condition_ready (fork15_outs_11_ready),
    .data (constant236_outs),
    .data_valid (constant236_outs_valid),
    .data_ready (constant236_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br67_trueOut),
    .trueOut_valid (cond_br67_trueOut_valid),
    .trueOut_ready (cond_br67_trueOut_ready),
    .falseOut (cond_br67_falseOut),
    .falseOut_valid (cond_br67_falseOut_valid),
    .falseOut_ready (cond_br67_falseOut_ready)
  );

  sink #(.DATA_TYPE(25)) sink55(
    .ins (cond_br67_falseOut),
    .ins_valid (cond_br67_falseOut_valid),
    .ins_ready (cond_br67_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(25), .OUTPUT_TYPE(27)) extsi120(
    .ins (cond_br67_trueOut),
    .ins_valid (cond_br67_trueOut_valid),
    .ins_ready (cond_br67_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi120_outs),
    .outs_valid (extsi120_outs_valid),
    .outs_ready (extsi120_outs_ready)
  );

  cond_br #(.DATA_TYPE(24)) cond_br68(
    .condition (fork15_outs_4),
    .condition_valid (fork15_outs_4_valid),
    .condition_ready (fork15_outs_4_ready),
    .data (constant147_outs),
    .data_valid (constant147_outs_valid),
    .data_ready (constant147_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br68_trueOut),
    .trueOut_valid (cond_br68_trueOut_valid),
    .trueOut_ready (cond_br68_trueOut_ready),
    .falseOut (cond_br68_falseOut),
    .falseOut_valid (cond_br68_falseOut_valid),
    .falseOut_ready (cond_br68_falseOut_ready)
  );

  sink #(.DATA_TYPE(24)) sink56(
    .ins (cond_br68_falseOut),
    .ins_valid (cond_br68_falseOut_valid),
    .ins_ready (cond_br68_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(16)) cond_br69(
    .condition (fork15_outs_10),
    .condition_valid (fork15_outs_10_valid),
    .condition_ready (fork15_outs_10_ready),
    .data (constant237_outs),
    .data_valid (constant237_outs_valid),
    .data_ready (constant237_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br69_trueOut),
    .trueOut_valid (cond_br69_trueOut_valid),
    .trueOut_ready (cond_br69_trueOut_ready),
    .falseOut (cond_br69_falseOut),
    .falseOut_valid (cond_br69_falseOut_valid),
    .falseOut_ready (cond_br69_falseOut_ready)
  );

  sink #(.DATA_TYPE(16)) sink57(
    .ins (cond_br69_falseOut),
    .ins_valid (cond_br69_falseOut_valid),
    .ins_ready (cond_br69_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(16), .OUTPUT_TYPE(21)) extsi121(
    .ins (cond_br69_trueOut),
    .ins_valid (cond_br69_trueOut_valid),
    .ins_ready (cond_br69_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi121_outs),
    .outs_valid (extsi121_outs_valid),
    .outs_ready (extsi121_outs_ready)
  );

  cond_br #(.DATA_TYPE(13)) cond_br70(
    .condition (fork15_outs_9),
    .condition_valid (fork15_outs_9_valid),
    .condition_ready (fork15_outs_9_ready),
    .data (constant238_outs),
    .data_valid (constant238_outs_valid),
    .data_ready (constant238_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br70_trueOut),
    .trueOut_valid (cond_br70_trueOut_valid),
    .trueOut_ready (cond_br70_trueOut_ready),
    .falseOut (cond_br70_falseOut),
    .falseOut_valid (cond_br70_falseOut_valid),
    .falseOut_ready (cond_br70_falseOut_ready)
  );

  sink #(.DATA_TYPE(13)) sink58(
    .ins (cond_br70_falseOut),
    .ins_valid (cond_br70_falseOut_valid),
    .ins_ready (cond_br70_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(13), .OUTPUT_TYPE(18)) extsi122(
    .ins (cond_br70_trueOut),
    .ins_valid (cond_br70_trueOut_valid),
    .ins_ready (cond_br70_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi122_outs),
    .outs_valid (extsi122_outs_valid),
    .outs_ready (extsi122_outs_ready)
  );

  cond_br #(.DATA_TYPE(14)) cond_br71(
    .condition (fork15_outs_3),
    .condition_valid (fork15_outs_3_valid),
    .condition_ready (fork15_outs_3_ready),
    .data (constant150_outs),
    .data_valid (constant150_outs_valid),
    .data_ready (constant150_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br71_trueOut),
    .trueOut_valid (cond_br71_trueOut_valid),
    .trueOut_ready (cond_br71_trueOut_ready),
    .falseOut (cond_br71_falseOut),
    .falseOut_valid (cond_br71_falseOut_valid),
    .falseOut_ready (cond_br71_falseOut_ready)
  );

  sink #(.DATA_TYPE(14)) sink59(
    .ins (cond_br71_falseOut),
    .ins_valid (cond_br71_falseOut_valid),
    .ins_ready (cond_br71_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br72(
    .condition (fork15_outs_2),
    .condition_valid (fork15_outs_2_valid),
    .condition_ready (fork15_outs_2_ready),
    .data (constant151_outs),
    .data_valid (constant151_outs_valid),
    .data_ready (constant151_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br72_trueOut),
    .trueOut_valid (cond_br72_trueOut_valid),
    .trueOut_ready (cond_br72_trueOut_ready),
    .falseOut (cond_br72_falseOut),
    .falseOut_valid (cond_br72_falseOut_valid),
    .falseOut_ready (cond_br72_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink60(
    .ins (cond_br72_falseOut),
    .ins_valid (cond_br72_falseOut_valid),
    .ins_ready (cond_br72_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(3)) cond_br73(
    .condition (fork15_outs_8),
    .condition_valid (fork15_outs_8_valid),
    .condition_ready (fork15_outs_8_ready),
    .data (constant234_outs),
    .data_valid (constant234_outs_valid),
    .data_ready (constant234_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br73_trueOut),
    .trueOut_valid (cond_br73_trueOut_valid),
    .trueOut_ready (cond_br73_trueOut_ready),
    .falseOut (cond_br73_falseOut),
    .falseOut_valid (cond_br73_falseOut_valid),
    .falseOut_ready (cond_br73_falseOut_ready)
  );

  sink #(.DATA_TYPE(3)) sink61(
    .ins (cond_br73_falseOut),
    .ins_valid (cond_br73_falseOut_valid),
    .ins_ready (cond_br73_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(8)) extsi123(
    .ins (cond_br73_trueOut),
    .ins_valid (cond_br73_trueOut_valid),
    .ins_ready (cond_br73_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi123_outs),
    .outs_valid (extsi123_outs_valid),
    .outs_ready (extsi123_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br74(
    .condition (fork15_outs_7),
    .condition_valid (fork15_outs_7_valid),
    .condition_ready (fork15_outs_7_ready),
    .data (constant239_outs),
    .data_valid (constant239_outs_valid),
    .data_ready (constant239_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br74_trueOut),
    .trueOut_valid (cond_br74_trueOut_valid),
    .trueOut_ready (cond_br74_trueOut_ready),
    .falseOut (cond_br74_falseOut),
    .falseOut_valid (cond_br74_falseOut_valid),
    .falseOut_ready (cond_br74_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink62(
    .ins (cond_br74_falseOut),
    .ins_valid (cond_br74_falseOut_valid),
    .ins_ready (cond_br74_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(8)) extsi124(
    .ins (cond_br74_trueOut),
    .ins_valid (cond_br74_trueOut_valid),
    .ins_ready (cond_br74_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi124_outs),
    .outs_valid (extsi124_outs_valid),
    .outs_ready (extsi124_outs_ready)
  );

  oehb #(.DATA_TYPE(5)) buffer18(
    .ins (cond_br61_falseOut),
    .ins_valid (cond_br61_falseOut_valid),
    .ins_ready (cond_br61_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer18_outs),
    .outs_valid (buffer18_outs_valid),
    .outs_ready (buffer18_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer19(
    .ins (buffer18_outs),
    .ins_valid (buffer18_outs_valid),
    .ins_ready (buffer18_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer19_outs),
    .outs_valid (buffer19_outs_valid),
    .outs_ready (buffer19_outs_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br75(
    .condition (fork15_outs_0),
    .condition_valid (fork15_outs_0_valid),
    .condition_ready (fork15_outs_0_ready),
    .data (buffer19_outs),
    .data_valid (buffer19_outs_valid),
    .data_ready (buffer19_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br75_trueOut),
    .trueOut_valid (cond_br75_trueOut_valid),
    .trueOut_ready (cond_br75_trueOut_ready),
    .falseOut (cond_br75_falseOut),
    .falseOut_valid (cond_br75_falseOut_valid),
    .falseOut_ready (cond_br75_falseOut_ready)
  );

  cond_br_dataless cond_br76(
    .condition (fork15_outs_1),
    .condition_valid (fork15_outs_1_valid),
    .condition_ready (fork15_outs_1_ready),
    .data_valid (fork14_outs_11_valid),
    .data_ready (fork14_outs_11_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br76_trueOut_valid),
    .trueOut_ready (cond_br76_trueOut_ready),
    .falseOut_valid (cond_br76_falseOut_valid),
    .falseOut_ready (cond_br76_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(3)) cond_br77(
    .condition (fork15_outs_13),
    .condition_valid (fork15_outs_13_valid),
    .condition_ready (fork15_outs_13_ready),
    .data (fork13_outs_1),
    .data_valid (fork13_outs_1_valid),
    .data_ready (fork13_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br77_trueOut),
    .trueOut_valid (cond_br77_trueOut_valid),
    .trueOut_ready (cond_br77_trueOut_ready),
    .falseOut (cond_br77_falseOut),
    .falseOut_valid (cond_br77_falseOut_valid),
    .falseOut_ready (cond_br77_falseOut_ready)
  );

  sink #(.DATA_TYPE(3)) sink63(
    .ins (cond_br77_trueOut),
    .ins_valid (cond_br77_trueOut_valid),
    .ins_ready (cond_br77_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(3)) buffer26(
    .ins (cond_br77_falseOut),
    .ins_valid (cond_br77_falseOut_valid),
    .ins_ready (cond_br77_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer26_outs),
    .outs_valid (buffer26_outs_valid),
    .outs_ready (buffer26_outs_ready)
  );

  tehb #(.DATA_TYPE(3)) buffer27(
    .ins (buffer26_outs),
    .ins_valid (buffer26_outs_valid),
    .ins_ready (buffer26_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer27_outs),
    .outs_valid (buffer27_outs_valid),
    .outs_ready (buffer27_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(3)) fork16(
    .ins (buffer27_outs),
    .ins_valid (buffer27_outs_valid),
    .ins_ready (buffer27_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork16_outs_1, fork16_outs_0}),
    .outs_valid ({fork16_outs_1_valid, fork16_outs_0_valid}),
    .outs_ready ({fork16_outs_1_ready, fork16_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(4)) extsi125(
    .ins (fork16_outs_0),
    .ins_valid (fork16_outs_0_valid),
    .ins_ready (fork16_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi125_outs),
    .outs_valid (extsi125_outs_valid),
    .outs_ready (extsi125_outs_ready)
  );

  oehb_dataless buffer28(
    .ins_valid (cond_br76_falseOut_valid),
    .ins_ready (cond_br76_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer28_outs_valid),
    .outs_ready (buffer28_outs_ready)
  );

  tehb_dataless buffer29(
    .ins_valid (buffer28_outs_valid),
    .ins_ready (buffer28_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer29_outs_valid),
    .outs_ready (buffer29_outs_ready)
  );

  fork_dataless #(.SIZE(12)) fork17(
    .ins_valid (buffer29_outs_valid),
    .ins_ready (buffer29_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork17_outs_11_valid, fork17_outs_10_valid, fork17_outs_9_valid, fork17_outs_8_valid, fork17_outs_7_valid, fork17_outs_6_valid, fork17_outs_5_valid, fork17_outs_4_valid, fork17_outs_3_valid, fork17_outs_2_valid, fork17_outs_1_valid, fork17_outs_0_valid}),
    .outs_ready ({fork17_outs_11_ready, fork17_outs_10_ready, fork17_outs_9_ready, fork17_outs_8_ready, fork17_outs_7_ready, fork17_outs_6_ready, fork17_outs_5_ready, fork17_outs_4_ready, fork17_outs_3_ready, fork17_outs_2_ready, fork17_outs_1_ready, fork17_outs_0_ready})
  );

  handshake_constant_1 #(.DATA_WIDTH(8)) constant154(
    .ctrl_valid (fork17_outs_10_valid),
    .ctrl_ready (fork17_outs_10_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant154_outs),
    .outs_valid (constant154_outs_valid),
    .outs_ready (constant154_outs_ready)
  );

  handshake_constant_59 #(.DATA_WIDTH(36)) constant155(
    .ctrl_valid (fork17_outs_9_valid),
    .ctrl_ready (fork17_outs_9_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant155_outs),
    .outs_valid (constant155_outs_valid),
    .outs_ready (constant155_outs_ready)
  );

  handshake_constant_60 #(.DATA_WIDTH(30)) constant241(
    .ctrl_valid (fork17_outs_4_valid),
    .ctrl_ready (fork17_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant241_outs),
    .outs_valid (constant241_outs_valid),
    .outs_ready (constant241_outs_ready)
  );

  handshake_constant_61 #(.DATA_WIDTH(30)) constant157(
    .ctrl_valid (fork17_outs_8_valid),
    .ctrl_ready (fork17_outs_8_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant157_outs),
    .outs_valid (constant157_outs_valid),
    .outs_ready (constant157_outs_ready)
  );

  handshake_constant_62 #(.DATA_WIDTH(24)) constant242(
    .ctrl_valid (fork17_outs_3_valid),
    .ctrl_ready (fork17_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant242_outs),
    .outs_valid (constant242_outs_valid),
    .outs_ready (constant242_outs_ready)
  );

  handshake_constant_63 #(.DATA_WIDTH(24)) constant159(
    .ctrl_valid (fork17_outs_7_valid),
    .ctrl_ready (fork17_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant159_outs),
    .outs_valid (constant159_outs_valid),
    .outs_ready (constant159_outs_ready)
  );

  handshake_constant_64 #(.DATA_WIDTH(17)) constant243(
    .ctrl_valid (fork17_outs_2_valid),
    .ctrl_ready (fork17_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant243_outs),
    .outs_valid (constant243_outs_valid),
    .outs_ready (constant243_outs_ready)
  );

  handshake_constant_65 #(.DATA_WIDTH(18)) constant161(
    .ctrl_valid (fork17_outs_6_valid),
    .ctrl_ready (fork17_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant161_outs),
    .outs_valid (constant161_outs_valid),
    .outs_ready (constant161_outs_ready)
  );

  handshake_constant_66 #(.DATA_WIDTH(14)) constant162(
    .ctrl_valid (fork17_outs_5_valid),
    .ctrl_ready (fork17_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant162_outs),
    .outs_valid (constant162_outs_valid),
    .outs_ready (constant162_outs_ready)
  );

  handshake_constant_67 #(.DATA_WIDTH(9)) constant244(
    .ctrl_valid (fork17_outs_1_valid),
    .ctrl_ready (fork17_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant244_outs),
    .outs_valid (constant244_outs_valid),
    .outs_ready (constant244_outs_ready)
  );

  handshake_constant_68 #(.DATA_WIDTH(6)) constant245(
    .ctrl_valid (fork17_outs_0_valid),
    .ctrl_ready (fork17_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant245_outs),
    .outs_valid (constant245_outs_valid),
    .outs_ready (constant245_outs_ready)
  );

  source source6(
    .clk (clk),
    .rst (rst),
    .outs_valid (source6_outs_valid),
    .outs_ready (source6_outs_ready)
  );

  handshake_constant_12 #(.DATA_WIDTH(4)) constant246(
    .ctrl_valid (source6_outs_valid),
    .ctrl_ready (source6_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant246_outs),
    .outs_valid (constant246_outs_valid),
    .outs_ready (constant246_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(4)) cmpi5(
    .lhs (extsi125_outs),
    .lhs_valid (extsi125_outs_valid),
    .lhs_ready (extsi125_outs_ready),
    .rhs (constant246_outs),
    .rhs_valid (constant246_outs_valid),
    .rhs_ready (constant246_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi5_result),
    .result_valid (cmpi5_result_valid),
    .result_ready (cmpi5_result_ready)
  );

  fork_type #(.SIZE(14), .DATA_TYPE(1)) fork18(
    .ins (cmpi5_result),
    .ins_valid (cmpi5_result_valid),
    .ins_ready (cmpi5_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork18_outs_13, fork18_outs_12, fork18_outs_11, fork18_outs_10, fork18_outs_9, fork18_outs_8, fork18_outs_7, fork18_outs_6, fork18_outs_5, fork18_outs_4, fork18_outs_3, fork18_outs_2, fork18_outs_1, fork18_outs_0}),
    .outs_valid ({fork18_outs_13_valid, fork18_outs_12_valid, fork18_outs_11_valid, fork18_outs_10_valid, fork18_outs_9_valid, fork18_outs_8_valid, fork18_outs_7_valid, fork18_outs_6_valid, fork18_outs_5_valid, fork18_outs_4_valid, fork18_outs_3_valid, fork18_outs_2_valid, fork18_outs_1_valid, fork18_outs_0_valid}),
    .outs_ready ({fork18_outs_13_ready, fork18_outs_12_ready, fork18_outs_11_ready, fork18_outs_10_ready, fork18_outs_9_ready, fork18_outs_8_ready, fork18_outs_7_ready, fork18_outs_6_ready, fork18_outs_5_ready, fork18_outs_4_ready, fork18_outs_3_ready, fork18_outs_2_ready, fork18_outs_1_ready, fork18_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(36)) cond_br78(
    .condition (fork18_outs_7),
    .condition_valid (fork18_outs_7_valid),
    .condition_ready (fork18_outs_7_ready),
    .data (constant155_outs),
    .data_valid (constant155_outs_valid),
    .data_ready (constant155_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br78_trueOut),
    .trueOut_valid (cond_br78_trueOut_valid),
    .trueOut_ready (cond_br78_trueOut_ready),
    .falseOut (cond_br78_falseOut),
    .falseOut_valid (cond_br78_falseOut_valid),
    .falseOut_ready (cond_br78_falseOut_ready)
  );

  sink #(.DATA_TYPE(36)) sink65(
    .ins (cond_br78_falseOut),
    .ins_valid (cond_br78_falseOut_valid),
    .ins_ready (cond_br78_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(30)) cond_br79(
    .condition (fork18_outs_12),
    .condition_valid (fork18_outs_12_valid),
    .condition_ready (fork18_outs_12_ready),
    .data (constant241_outs),
    .data_valid (constant241_outs_valid),
    .data_ready (constant241_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br79_trueOut),
    .trueOut_valid (cond_br79_trueOut_valid),
    .trueOut_ready (cond_br79_trueOut_ready),
    .falseOut (cond_br79_falseOut),
    .falseOut_valid (cond_br79_falseOut_valid),
    .falseOut_ready (cond_br79_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink66(
    .ins (cond_br79_falseOut),
    .ins_valid (cond_br79_falseOut_valid),
    .ins_ready (cond_br79_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(30), .OUTPUT_TYPE(34)) extsi126(
    .ins (cond_br79_trueOut),
    .ins_valid (cond_br79_trueOut_valid),
    .ins_ready (cond_br79_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi126_outs),
    .outs_valid (extsi126_outs_valid),
    .outs_ready (extsi126_outs_ready)
  );

  cond_br #(.DATA_TYPE(30)) cond_br80(
    .condition (fork18_outs_6),
    .condition_valid (fork18_outs_6_valid),
    .condition_ready (fork18_outs_6_ready),
    .data (constant157_outs),
    .data_valid (constant157_outs_valid),
    .data_ready (constant157_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br80_trueOut),
    .trueOut_valid (cond_br80_trueOut_valid),
    .trueOut_ready (cond_br80_trueOut_ready),
    .falseOut (cond_br80_falseOut),
    .falseOut_valid (cond_br80_falseOut_valid),
    .falseOut_ready (cond_br80_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink67(
    .ins (cond_br80_falseOut),
    .ins_valid (cond_br80_falseOut_valid),
    .ins_ready (cond_br80_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(24)) cond_br81(
    .condition (fork18_outs_11),
    .condition_valid (fork18_outs_11_valid),
    .condition_ready (fork18_outs_11_ready),
    .data (constant242_outs),
    .data_valid (constant242_outs_valid),
    .data_ready (constant242_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br81_trueOut),
    .trueOut_valid (cond_br81_trueOut_valid),
    .trueOut_ready (cond_br81_trueOut_ready),
    .falseOut (cond_br81_falseOut),
    .falseOut_valid (cond_br81_falseOut_valid),
    .falseOut_ready (cond_br81_falseOut_ready)
  );

  sink #(.DATA_TYPE(24)) sink68(
    .ins (cond_br81_falseOut),
    .ins_valid (cond_br81_falseOut_valid),
    .ins_ready (cond_br81_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(24), .OUTPUT_TYPE(27)) extsi127(
    .ins (cond_br81_trueOut),
    .ins_valid (cond_br81_trueOut_valid),
    .ins_ready (cond_br81_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi127_outs),
    .outs_valid (extsi127_outs_valid),
    .outs_ready (extsi127_outs_ready)
  );

  cond_br #(.DATA_TYPE(24)) cond_br82(
    .condition (fork18_outs_5),
    .condition_valid (fork18_outs_5_valid),
    .condition_ready (fork18_outs_5_ready),
    .data (constant159_outs),
    .data_valid (constant159_outs_valid),
    .data_ready (constant159_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br82_trueOut),
    .trueOut_valid (cond_br82_trueOut_valid),
    .trueOut_ready (cond_br82_trueOut_ready),
    .falseOut (cond_br82_falseOut),
    .falseOut_valid (cond_br82_falseOut_valid),
    .falseOut_ready (cond_br82_falseOut_ready)
  );

  sink #(.DATA_TYPE(24)) sink69(
    .ins (cond_br82_falseOut),
    .ins_valid (cond_br82_falseOut_valid),
    .ins_ready (cond_br82_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(17)) cond_br83(
    .condition (fork18_outs_10),
    .condition_valid (fork18_outs_10_valid),
    .condition_ready (fork18_outs_10_ready),
    .data (constant243_outs),
    .data_valid (constant243_outs_valid),
    .data_ready (constant243_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br83_trueOut),
    .trueOut_valid (cond_br83_trueOut_valid),
    .trueOut_ready (cond_br83_trueOut_ready),
    .falseOut (cond_br83_falseOut),
    .falseOut_valid (cond_br83_falseOut_valid),
    .falseOut_ready (cond_br83_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink70(
    .ins (cond_br83_falseOut),
    .ins_valid (cond_br83_falseOut_valid),
    .ins_ready (cond_br83_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(17), .OUTPUT_TYPE(21)) extsi128(
    .ins (cond_br83_trueOut),
    .ins_valid (cond_br83_trueOut_valid),
    .ins_ready (cond_br83_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi128_outs),
    .outs_valid (extsi128_outs_valid),
    .outs_ready (extsi128_outs_ready)
  );

  cond_br #(.DATA_TYPE(18)) cond_br84(
    .condition (fork18_outs_4),
    .condition_valid (fork18_outs_4_valid),
    .condition_ready (fork18_outs_4_ready),
    .data (constant161_outs),
    .data_valid (constant161_outs_valid),
    .data_ready (constant161_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br84_trueOut),
    .trueOut_valid (cond_br84_trueOut_valid),
    .trueOut_ready (cond_br84_trueOut_ready),
    .falseOut (cond_br84_falseOut),
    .falseOut_valid (cond_br84_falseOut_valid),
    .falseOut_ready (cond_br84_falseOut_ready)
  );

  sink #(.DATA_TYPE(18)) sink71(
    .ins (cond_br84_falseOut),
    .ins_valid (cond_br84_falseOut_valid),
    .ins_ready (cond_br84_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(14)) cond_br85(
    .condition (fork18_outs_3),
    .condition_valid (fork18_outs_3_valid),
    .condition_ready (fork18_outs_3_ready),
    .data (constant162_outs),
    .data_valid (constant162_outs_valid),
    .data_ready (constant162_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br85_trueOut),
    .trueOut_valid (cond_br85_trueOut_valid),
    .trueOut_ready (cond_br85_trueOut_ready),
    .falseOut (cond_br85_falseOut),
    .falseOut_valid (cond_br85_falseOut_valid),
    .falseOut_ready (cond_br85_falseOut_ready)
  );

  sink #(.DATA_TYPE(14)) sink72(
    .ins (cond_br85_falseOut),
    .ins_valid (cond_br85_falseOut_valid),
    .ins_ready (cond_br85_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(9)) cond_br86(
    .condition (fork18_outs_9),
    .condition_valid (fork18_outs_9_valid),
    .condition_ready (fork18_outs_9_ready),
    .data (constant244_outs),
    .data_valid (constant244_outs_valid),
    .data_ready (constant244_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br86_trueOut),
    .trueOut_valid (cond_br86_trueOut_valid),
    .trueOut_ready (cond_br86_trueOut_ready),
    .falseOut (cond_br86_falseOut),
    .falseOut_valid (cond_br86_falseOut_valid),
    .falseOut_ready (cond_br86_falseOut_ready)
  );

  sink #(.DATA_TYPE(9)) sink73(
    .ins (cond_br86_falseOut),
    .ins_valid (cond_br86_falseOut_valid),
    .ins_ready (cond_br86_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(9), .OUTPUT_TYPE(12)) extsi129(
    .ins (cond_br86_trueOut),
    .ins_valid (cond_br86_trueOut_valid),
    .ins_ready (cond_br86_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi129_outs),
    .outs_valid (extsi129_outs_valid),
    .outs_ready (extsi129_outs_ready)
  );

  cond_br #(.DATA_TYPE(6)) cond_br87(
    .condition (fork18_outs_8),
    .condition_valid (fork18_outs_8_valid),
    .condition_ready (fork18_outs_8_ready),
    .data (constant245_outs),
    .data_valid (constant245_outs_valid),
    .data_ready (constant245_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br87_trueOut),
    .trueOut_valid (cond_br87_trueOut_valid),
    .trueOut_ready (cond_br87_trueOut_ready),
    .falseOut (cond_br87_falseOut),
    .falseOut_valid (cond_br87_falseOut_valid),
    .falseOut_ready (cond_br87_falseOut_ready)
  );

  sink #(.DATA_TYPE(6)) sink74(
    .ins (cond_br87_falseOut),
    .ins_valid (cond_br87_falseOut_valid),
    .ins_ready (cond_br87_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(8)) extsi130(
    .ins (cond_br87_trueOut),
    .ins_valid (cond_br87_trueOut_valid),
    .ins_ready (cond_br87_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi130_outs),
    .outs_valid (extsi130_outs_valid),
    .outs_ready (extsi130_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br88(
    .condition (fork18_outs_2),
    .condition_valid (fork18_outs_2_valid),
    .condition_ready (fork18_outs_2_ready),
    .data (constant154_outs),
    .data_valid (constant154_outs_valid),
    .data_ready (constant154_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br88_trueOut),
    .trueOut_valid (cond_br88_trueOut_valid),
    .trueOut_ready (cond_br88_trueOut_ready),
    .falseOut (cond_br88_falseOut),
    .falseOut_valid (cond_br88_falseOut_valid),
    .falseOut_ready (cond_br88_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink75(
    .ins (cond_br88_falseOut),
    .ins_valid (cond_br88_falseOut_valid),
    .ins_ready (cond_br88_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer24(
    .ins (cond_br75_falseOut),
    .ins_valid (cond_br75_falseOut_valid),
    .ins_ready (cond_br75_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer24_outs),
    .outs_valid (buffer24_outs_valid),
    .outs_ready (buffer24_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer25(
    .ins (buffer24_outs),
    .ins_valid (buffer24_outs_valid),
    .ins_ready (buffer24_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer25_outs),
    .outs_valid (buffer25_outs_valid),
    .outs_ready (buffer25_outs_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br89(
    .condition (fork18_outs_0),
    .condition_valid (fork18_outs_0_valid),
    .condition_ready (fork18_outs_0_ready),
    .data (buffer25_outs),
    .data_valid (buffer25_outs_valid),
    .data_ready (buffer25_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br89_trueOut),
    .trueOut_valid (cond_br89_trueOut_valid),
    .trueOut_ready (cond_br89_trueOut_ready),
    .falseOut (cond_br89_falseOut),
    .falseOut_valid (cond_br89_falseOut_valid),
    .falseOut_ready (cond_br89_falseOut_ready)
  );

  cond_br_dataless cond_br90(
    .condition (fork18_outs_1),
    .condition_valid (fork18_outs_1_valid),
    .condition_ready (fork18_outs_1_ready),
    .data_valid (fork17_outs_11_valid),
    .data_ready (fork17_outs_11_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br90_trueOut_valid),
    .trueOut_ready (cond_br90_trueOut_ready),
    .falseOut_valid (cond_br90_falseOut_valid),
    .falseOut_ready (cond_br90_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(3)) cond_br91(
    .condition (fork18_outs_13),
    .condition_valid (fork18_outs_13_valid),
    .condition_ready (fork18_outs_13_ready),
    .data (fork16_outs_1),
    .data_valid (fork16_outs_1_valid),
    .data_ready (fork16_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br91_trueOut),
    .trueOut_valid (cond_br91_trueOut_valid),
    .trueOut_ready (cond_br91_trueOut_ready),
    .falseOut (cond_br91_falseOut),
    .falseOut_valid (cond_br91_falseOut_valid),
    .falseOut_ready (cond_br91_falseOut_ready)
  );

  sink #(.DATA_TYPE(3)) sink76(
    .ins (cond_br91_trueOut),
    .ins_valid (cond_br91_trueOut_valid),
    .ins_ready (cond_br91_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(3)) buffer32(
    .ins (cond_br91_falseOut),
    .ins_valid (cond_br91_falseOut_valid),
    .ins_ready (cond_br91_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer32_outs),
    .outs_valid (buffer32_outs_valid),
    .outs_ready (buffer32_outs_ready)
  );

  tehb #(.DATA_TYPE(3)) buffer33(
    .ins (buffer32_outs),
    .ins_valid (buffer32_outs_valid),
    .ins_ready (buffer32_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer33_outs),
    .outs_valid (buffer33_outs_valid),
    .outs_ready (buffer33_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(3)) fork19(
    .ins (buffer33_outs),
    .ins_valid (buffer33_outs_valid),
    .ins_ready (buffer33_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork19_outs_1, fork19_outs_0}),
    .outs_valid ({fork19_outs_1_valid, fork19_outs_0_valid}),
    .outs_ready ({fork19_outs_1_ready, fork19_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(4)) extsi131(
    .ins (fork19_outs_0),
    .ins_valid (fork19_outs_0_valid),
    .ins_ready (fork19_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi131_outs),
    .outs_valid (extsi131_outs_valid),
    .outs_ready (extsi131_outs_ready)
  );

  oehb_dataless buffer34(
    .ins_valid (cond_br90_falseOut_valid),
    .ins_ready (cond_br90_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer34_outs_valid),
    .outs_ready (buffer34_outs_ready)
  );

  tehb_dataless buffer35(
    .ins_valid (buffer34_outs_valid),
    .ins_ready (buffer34_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer35_outs_valid),
    .outs_ready (buffer35_outs_ready)
  );

  fork_dataless #(.SIZE(12)) fork20(
    .ins_valid (buffer35_outs_valid),
    .ins_ready (buffer35_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork20_outs_11_valid, fork20_outs_10_valid, fork20_outs_9_valid, fork20_outs_8_valid, fork20_outs_7_valid, fork20_outs_6_valid, fork20_outs_5_valid, fork20_outs_4_valid, fork20_outs_3_valid, fork20_outs_2_valid, fork20_outs_1_valid, fork20_outs_0_valid}),
    .outs_ready ({fork20_outs_11_ready, fork20_outs_10_ready, fork20_outs_9_ready, fork20_outs_8_ready, fork20_outs_7_ready, fork20_outs_6_ready, fork20_outs_5_ready, fork20_outs_4_ready, fork20_outs_3_ready, fork20_outs_2_ready, fork20_outs_1_ready, fork20_outs_0_ready})
  );

  handshake_constant_69 #(.DATA_WIDTH(36)) constant166(
    .ctrl_valid (fork20_outs_10_valid),
    .ctrl_ready (fork20_outs_10_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant166_outs),
    .outs_valid (constant166_outs_valid),
    .outs_ready (constant166_outs_ready)
  );

  handshake_constant_70 #(.DATA_WIDTH(29)) constant247(
    .ctrl_valid (fork20_outs_4_valid),
    .ctrl_ready (fork20_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant247_outs),
    .outs_valid (constant247_outs_valid),
    .outs_ready (constant247_outs_ready)
  );

  handshake_constant_71 #(.DATA_WIDTH(30)) constant168(
    .ctrl_valid (fork20_outs_9_valid),
    .ctrl_ready (fork20_outs_9_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant168_outs),
    .outs_valid (constant168_outs_valid),
    .outs_ready (constant168_outs_ready)
  );

  handshake_constant_72 #(.DATA_WIDTH(23)) constant248(
    .ctrl_valid (fork20_outs_3_valid),
    .ctrl_ready (fork20_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant248_outs),
    .outs_valid (constant248_outs_valid),
    .outs_ready (constant248_outs_ready)
  );

  handshake_constant_73 #(.DATA_WIDTH(24)) constant170(
    .ctrl_valid (fork20_outs_8_valid),
    .ctrl_ready (fork20_outs_8_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant170_outs),
    .outs_valid (constant170_outs_valid),
    .outs_ready (constant170_outs_ready)
  );

  handshake_constant_74 #(.DATA_WIDTH(16)) constant249(
    .ctrl_valid (fork20_outs_2_valid),
    .ctrl_ready (fork20_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant249_outs),
    .outs_valid (constant249_outs_valid),
    .outs_ready (constant249_outs_ready)
  );

  handshake_constant_75 #(.DATA_WIDTH(18)) constant172(
    .ctrl_valid (fork20_outs_7_valid),
    .ctrl_ready (fork20_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant172_outs),
    .outs_valid (constant172_outs_valid),
    .outs_ready (constant172_outs_ready)
  );

  handshake_constant_68 #(.DATA_WIDTH(6)) constant250(
    .ctrl_valid (fork20_outs_1_valid),
    .ctrl_ready (fork20_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant250_outs),
    .outs_valid (constant250_outs_valid),
    .outs_ready (constant250_outs_ready)
  );

  handshake_constant_76 #(.DATA_WIDTH(12)) constant174(
    .ctrl_valid (fork20_outs_6_valid),
    .ctrl_ready (fork20_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant174_outs),
    .outs_valid (constant174_outs_valid),
    .outs_ready (constant174_outs_ready)
  );

  handshake_constant_77 #(.DATA_WIDTH(8)) constant175(
    .ctrl_valid (fork20_outs_5_valid),
    .ctrl_ready (fork20_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant175_outs),
    .outs_valid (constant175_outs_valid),
    .outs_ready (constant175_outs_ready)
  );

  handshake_constant_78 #(.DATA_WIDTH(5)) constant251(
    .ctrl_valid (fork20_outs_0_valid),
    .ctrl_ready (fork20_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant251_outs),
    .outs_valid (constant251_outs_valid),
    .outs_ready (constant251_outs_ready)
  );

  source source7(
    .clk (clk),
    .rst (rst),
    .outs_valid (source7_outs_valid),
    .outs_ready (source7_outs_ready)
  );

  handshake_constant_79 #(.DATA_WIDTH(4)) constant252(
    .ctrl_valid (source7_outs_valid),
    .ctrl_ready (source7_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant252_outs),
    .outs_valid (constant252_outs_valid),
    .outs_ready (constant252_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(4)) cmpi6(
    .lhs (extsi131_outs),
    .lhs_valid (extsi131_outs_valid),
    .lhs_ready (extsi131_outs_ready),
    .rhs (constant252_outs),
    .rhs_valid (constant252_outs_valid),
    .rhs_ready (constant252_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi6_result),
    .result_valid (cmpi6_result_valid),
    .result_ready (cmpi6_result_ready)
  );

  fork_type #(.SIZE(14), .DATA_TYPE(1)) fork21(
    .ins (cmpi6_result),
    .ins_valid (cmpi6_result_valid),
    .ins_ready (cmpi6_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork21_outs_13, fork21_outs_12, fork21_outs_11, fork21_outs_10, fork21_outs_9, fork21_outs_8, fork21_outs_7, fork21_outs_6, fork21_outs_5, fork21_outs_4, fork21_outs_3, fork21_outs_2, fork21_outs_1, fork21_outs_0}),
    .outs_valid ({fork21_outs_13_valid, fork21_outs_12_valid, fork21_outs_11_valid, fork21_outs_10_valid, fork21_outs_9_valid, fork21_outs_8_valid, fork21_outs_7_valid, fork21_outs_6_valid, fork21_outs_5_valid, fork21_outs_4_valid, fork21_outs_3_valid, fork21_outs_2_valid, fork21_outs_1_valid, fork21_outs_0_valid}),
    .outs_ready ({fork21_outs_13_ready, fork21_outs_12_ready, fork21_outs_11_ready, fork21_outs_10_ready, fork21_outs_9_ready, fork21_outs_8_ready, fork21_outs_7_ready, fork21_outs_6_ready, fork21_outs_5_ready, fork21_outs_4_ready, fork21_outs_3_ready, fork21_outs_2_ready, fork21_outs_1_ready, fork21_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(36)) cond_br92(
    .condition (fork21_outs_7),
    .condition_valid (fork21_outs_7_valid),
    .condition_ready (fork21_outs_7_ready),
    .data (constant166_outs),
    .data_valid (constant166_outs_valid),
    .data_ready (constant166_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br92_trueOut),
    .trueOut_valid (cond_br92_trueOut_valid),
    .trueOut_ready (cond_br92_trueOut_ready),
    .falseOut (cond_br92_falseOut),
    .falseOut_valid (cond_br92_falseOut_valid),
    .falseOut_ready (cond_br92_falseOut_ready)
  );

  sink #(.DATA_TYPE(36)) sink78(
    .ins (cond_br92_falseOut),
    .ins_valid (cond_br92_falseOut_valid),
    .ins_ready (cond_br92_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(29)) cond_br93(
    .condition (fork21_outs_12),
    .condition_valid (fork21_outs_12_valid),
    .condition_ready (fork21_outs_12_ready),
    .data (constant247_outs),
    .data_valid (constant247_outs_valid),
    .data_ready (constant247_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br93_trueOut),
    .trueOut_valid (cond_br93_trueOut_valid),
    .trueOut_ready (cond_br93_trueOut_ready),
    .falseOut (cond_br93_falseOut),
    .falseOut_valid (cond_br93_falseOut_valid),
    .falseOut_ready (cond_br93_falseOut_ready)
  );

  sink #(.DATA_TYPE(29)) sink79(
    .ins (cond_br93_falseOut),
    .ins_valid (cond_br93_falseOut_valid),
    .ins_ready (cond_br93_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(29), .OUTPUT_TYPE(34)) extsi132(
    .ins (cond_br93_trueOut),
    .ins_valid (cond_br93_trueOut_valid),
    .ins_ready (cond_br93_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi132_outs),
    .outs_valid (extsi132_outs_valid),
    .outs_ready (extsi132_outs_ready)
  );

  cond_br #(.DATA_TYPE(30)) cond_br94(
    .condition (fork21_outs_6),
    .condition_valid (fork21_outs_6_valid),
    .condition_ready (fork21_outs_6_ready),
    .data (constant168_outs),
    .data_valid (constant168_outs_valid),
    .data_ready (constant168_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br94_trueOut),
    .trueOut_valid (cond_br94_trueOut_valid),
    .trueOut_ready (cond_br94_trueOut_ready),
    .falseOut (cond_br94_falseOut),
    .falseOut_valid (cond_br94_falseOut_valid),
    .falseOut_ready (cond_br94_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink80(
    .ins (cond_br94_falseOut),
    .ins_valid (cond_br94_falseOut_valid),
    .ins_ready (cond_br94_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(23)) cond_br95(
    .condition (fork21_outs_11),
    .condition_valid (fork21_outs_11_valid),
    .condition_ready (fork21_outs_11_ready),
    .data (constant248_outs),
    .data_valid (constant248_outs_valid),
    .data_ready (constant248_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br95_trueOut),
    .trueOut_valid (cond_br95_trueOut_valid),
    .trueOut_ready (cond_br95_trueOut_ready),
    .falseOut (cond_br95_falseOut),
    .falseOut_valid (cond_br95_falseOut_valid),
    .falseOut_ready (cond_br95_falseOut_ready)
  );

  sink #(.DATA_TYPE(23)) sink81(
    .ins (cond_br95_falseOut),
    .ins_valid (cond_br95_falseOut_valid),
    .ins_ready (cond_br95_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(23), .OUTPUT_TYPE(27)) extsi133(
    .ins (cond_br95_trueOut),
    .ins_valid (cond_br95_trueOut_valid),
    .ins_ready (cond_br95_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi133_outs),
    .outs_valid (extsi133_outs_valid),
    .outs_ready (extsi133_outs_ready)
  );

  cond_br #(.DATA_TYPE(24)) cond_br96(
    .condition (fork21_outs_5),
    .condition_valid (fork21_outs_5_valid),
    .condition_ready (fork21_outs_5_ready),
    .data (constant170_outs),
    .data_valid (constant170_outs_valid),
    .data_ready (constant170_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br96_trueOut),
    .trueOut_valid (cond_br96_trueOut_valid),
    .trueOut_ready (cond_br96_trueOut_ready),
    .falseOut (cond_br96_falseOut),
    .falseOut_valid (cond_br96_falseOut_valid),
    .falseOut_ready (cond_br96_falseOut_ready)
  );

  sink #(.DATA_TYPE(24)) sink82(
    .ins (cond_br96_falseOut),
    .ins_valid (cond_br96_falseOut_valid),
    .ins_ready (cond_br96_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(16)) cond_br97(
    .condition (fork21_outs_10),
    .condition_valid (fork21_outs_10_valid),
    .condition_ready (fork21_outs_10_ready),
    .data (constant249_outs),
    .data_valid (constant249_outs_valid),
    .data_ready (constant249_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br97_trueOut),
    .trueOut_valid (cond_br97_trueOut_valid),
    .trueOut_ready (cond_br97_trueOut_ready),
    .falseOut (cond_br97_falseOut),
    .falseOut_valid (cond_br97_falseOut_valid),
    .falseOut_ready (cond_br97_falseOut_ready)
  );

  sink #(.DATA_TYPE(16)) sink83(
    .ins (cond_br97_falseOut),
    .ins_valid (cond_br97_falseOut_valid),
    .ins_ready (cond_br97_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(16), .OUTPUT_TYPE(21)) extsi134(
    .ins (cond_br97_trueOut),
    .ins_valid (cond_br97_trueOut_valid),
    .ins_ready (cond_br97_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi134_outs),
    .outs_valid (extsi134_outs_valid),
    .outs_ready (extsi134_outs_ready)
  );

  cond_br #(.DATA_TYPE(18)) cond_br98(
    .condition (fork21_outs_4),
    .condition_valid (fork21_outs_4_valid),
    .condition_ready (fork21_outs_4_ready),
    .data (constant172_outs),
    .data_valid (constant172_outs_valid),
    .data_ready (constant172_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br98_trueOut),
    .trueOut_valid (cond_br98_trueOut_valid),
    .trueOut_ready (cond_br98_trueOut_ready),
    .falseOut (cond_br98_falseOut),
    .falseOut_valid (cond_br98_falseOut_valid),
    .falseOut_ready (cond_br98_falseOut_ready)
  );

  sink #(.DATA_TYPE(18)) sink84(
    .ins (cond_br98_falseOut),
    .ins_valid (cond_br98_falseOut_valid),
    .ins_ready (cond_br98_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(6)) cond_br99(
    .condition (fork21_outs_9),
    .condition_valid (fork21_outs_9_valid),
    .condition_ready (fork21_outs_9_ready),
    .data (constant250_outs),
    .data_valid (constant250_outs_valid),
    .data_ready (constant250_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br99_trueOut),
    .trueOut_valid (cond_br99_trueOut_valid),
    .trueOut_ready (cond_br99_trueOut_ready),
    .falseOut (cond_br99_falseOut),
    .falseOut_valid (cond_br99_falseOut_valid),
    .falseOut_ready (cond_br99_falseOut_ready)
  );

  sink #(.DATA_TYPE(6)) sink85(
    .ins (cond_br99_falseOut),
    .ins_valid (cond_br99_falseOut_valid),
    .ins_ready (cond_br99_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(14)) extsi135(
    .ins (cond_br99_trueOut),
    .ins_valid (cond_br99_trueOut_valid),
    .ins_ready (cond_br99_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi135_outs),
    .outs_valid (extsi135_outs_valid),
    .outs_ready (extsi135_outs_ready)
  );

  cond_br #(.DATA_TYPE(12)) cond_br100(
    .condition (fork21_outs_3),
    .condition_valid (fork21_outs_3_valid),
    .condition_ready (fork21_outs_3_ready),
    .data (constant174_outs),
    .data_valid (constant174_outs_valid),
    .data_ready (constant174_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br100_trueOut),
    .trueOut_valid (cond_br100_trueOut_valid),
    .trueOut_ready (cond_br100_trueOut_ready),
    .falseOut (cond_br100_falseOut),
    .falseOut_valid (cond_br100_falseOut_valid),
    .falseOut_ready (cond_br100_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink86(
    .ins (cond_br100_falseOut),
    .ins_valid (cond_br100_falseOut_valid),
    .ins_ready (cond_br100_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(8)) cond_br101(
    .condition (fork21_outs_2),
    .condition_valid (fork21_outs_2_valid),
    .condition_ready (fork21_outs_2_ready),
    .data (constant175_outs),
    .data_valid (constant175_outs_valid),
    .data_ready (constant175_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br101_trueOut),
    .trueOut_valid (cond_br101_trueOut_valid),
    .trueOut_ready (cond_br101_trueOut_ready),
    .falseOut (cond_br101_falseOut),
    .falseOut_valid (cond_br101_falseOut_valid),
    .falseOut_ready (cond_br101_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink87(
    .ins (cond_br101_falseOut),
    .ins_valid (cond_br101_falseOut_valid),
    .ins_ready (cond_br101_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(5)) cond_br102(
    .condition (fork21_outs_8),
    .condition_valid (fork21_outs_8_valid),
    .condition_ready (fork21_outs_8_ready),
    .data (constant251_outs),
    .data_valid (constant251_outs_valid),
    .data_ready (constant251_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br102_trueOut),
    .trueOut_valid (cond_br102_trueOut_valid),
    .trueOut_ready (cond_br102_trueOut_ready),
    .falseOut (cond_br102_falseOut),
    .falseOut_valid (cond_br102_falseOut_valid),
    .falseOut_ready (cond_br102_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink88(
    .ins (cond_br102_falseOut),
    .ins_valid (cond_br102_falseOut_valid),
    .ins_ready (cond_br102_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(8)) extsi136(
    .ins (cond_br102_trueOut),
    .ins_valid (cond_br102_trueOut_valid),
    .ins_ready (cond_br102_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi136_outs),
    .outs_valid (extsi136_outs_valid),
    .outs_ready (extsi136_outs_ready)
  );

  oehb #(.DATA_TYPE(5)) buffer30(
    .ins (cond_br89_falseOut),
    .ins_valid (cond_br89_falseOut_valid),
    .ins_ready (cond_br89_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer30_outs),
    .outs_valid (buffer30_outs_valid),
    .outs_ready (buffer30_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer31(
    .ins (buffer30_outs),
    .ins_valid (buffer30_outs_valid),
    .ins_ready (buffer30_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer31_outs),
    .outs_valid (buffer31_outs_valid),
    .outs_ready (buffer31_outs_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br103(
    .condition (fork21_outs_0),
    .condition_valid (fork21_outs_0_valid),
    .condition_ready (fork21_outs_0_ready),
    .data (buffer31_outs),
    .data_valid (buffer31_outs_valid),
    .data_ready (buffer31_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br103_trueOut),
    .trueOut_valid (cond_br103_trueOut_valid),
    .trueOut_ready (cond_br103_trueOut_ready),
    .falseOut (cond_br103_falseOut),
    .falseOut_valid (cond_br103_falseOut_valid),
    .falseOut_ready (cond_br103_falseOut_ready)
  );

  cond_br_dataless cond_br104(
    .condition (fork21_outs_1),
    .condition_valid (fork21_outs_1_valid),
    .condition_ready (fork21_outs_1_ready),
    .data_valid (fork20_outs_11_valid),
    .data_ready (fork20_outs_11_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br104_trueOut_valid),
    .trueOut_ready (cond_br104_trueOut_ready),
    .falseOut_valid (cond_br104_falseOut_valid),
    .falseOut_ready (cond_br104_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(3)) cond_br105(
    .condition (fork21_outs_13),
    .condition_valid (fork21_outs_13_valid),
    .condition_ready (fork21_outs_13_ready),
    .data (fork19_outs_1),
    .data_valid (fork19_outs_1_valid),
    .data_ready (fork19_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br105_trueOut),
    .trueOut_valid (cond_br105_trueOut_valid),
    .trueOut_ready (cond_br105_trueOut_ready),
    .falseOut (cond_br105_falseOut),
    .falseOut_valid (cond_br105_falseOut_valid),
    .falseOut_ready (cond_br105_falseOut_ready)
  );

  sink #(.DATA_TYPE(3)) sink89(
    .ins (cond_br105_trueOut),
    .ins_valid (cond_br105_trueOut_valid),
    .ins_ready (cond_br105_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(3)) buffer38(
    .ins (cond_br105_falseOut),
    .ins_valid (cond_br105_falseOut_valid),
    .ins_ready (cond_br105_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer38_outs),
    .outs_valid (buffer38_outs_valid),
    .outs_ready (buffer38_outs_ready)
  );

  tehb #(.DATA_TYPE(3)) buffer39(
    .ins (buffer38_outs),
    .ins_valid (buffer38_outs_valid),
    .ins_ready (buffer38_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer39_outs),
    .outs_valid (buffer39_outs_valid),
    .outs_ready (buffer39_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(4)) extsi137(
    .ins (buffer39_outs),
    .ins_valid (buffer39_outs_valid),
    .ins_ready (buffer39_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi137_outs),
    .outs_valid (extsi137_outs_valid),
    .outs_ready (extsi137_outs_ready)
  );

  oehb_dataless buffer40(
    .ins_valid (cond_br104_falseOut_valid),
    .ins_ready (cond_br104_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer40_outs_valid),
    .outs_ready (buffer40_outs_ready)
  );

  tehb_dataless buffer41(
    .ins_valid (buffer40_outs_valid),
    .ins_ready (buffer40_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer41_outs_valid),
    .outs_ready (buffer41_outs_ready)
  );

  fork_dataless #(.SIZE(23)) fork22(
    .ins_valid (buffer41_outs_valid),
    .ins_ready (buffer41_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork22_outs_22_valid, fork22_outs_21_valid, fork22_outs_20_valid, fork22_outs_19_valid, fork22_outs_18_valid, fork22_outs_17_valid, fork22_outs_16_valid, fork22_outs_15_valid, fork22_outs_14_valid, fork22_outs_13_valid, fork22_outs_12_valid, fork22_outs_11_valid, fork22_outs_10_valid, fork22_outs_9_valid, fork22_outs_8_valid, fork22_outs_7_valid, fork22_outs_6_valid, fork22_outs_5_valid, fork22_outs_4_valid, fork22_outs_3_valid, fork22_outs_2_valid, fork22_outs_1_valid, fork22_outs_0_valid}),
    .outs_ready ({fork22_outs_22_ready, fork22_outs_21_ready, fork22_outs_20_ready, fork22_outs_19_ready, fork22_outs_18_ready, fork22_outs_17_ready, fork22_outs_16_ready, fork22_outs_15_ready, fork22_outs_14_ready, fork22_outs_13_ready, fork22_outs_12_ready, fork22_outs_11_ready, fork22_outs_10_ready, fork22_outs_9_ready, fork22_outs_8_ready, fork22_outs_7_ready, fork22_outs_6_ready, fork22_outs_5_ready, fork22_outs_4_ready, fork22_outs_3_ready, fork22_outs_2_ready, fork22_outs_1_ready, fork22_outs_0_ready})
  );

  handshake_constant_11 #(.DATA_WIDTH(34)) constant253(
    .ctrl_valid (fork22_outs_5_valid),
    .ctrl_ready (fork22_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant253_outs),
    .outs_valid (constant253_outs_valid),
    .outs_ready (constant253_outs_ready)
  );

  handshake_constant_10 #(.DATA_WIDTH(34)) constant179(
    .ctrl_valid (fork22_outs_21_valid),
    .ctrl_ready (fork22_outs_21_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant179_outs),
    .outs_valid (constant179_outs_valid),
    .outs_ready (constant179_outs_ready)
  );

  handshake_constant_9 #(.DATA_WIDTH(30)) constant180(
    .ctrl_valid (fork22_outs_20_valid),
    .ctrl_ready (fork22_outs_20_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant180_outs),
    .outs_valid (constant180_outs_valid),
    .outs_ready (constant180_outs_ready)
  );

  handshake_constant_8 #(.DATA_WIDTH(27)) constant181(
    .ctrl_valid (fork22_outs_19_valid),
    .ctrl_ready (fork22_outs_19_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant181_outs),
    .outs_valid (constant181_outs_valid),
    .outs_ready (constant181_outs_ready)
  );

  handshake_constant_7 #(.DATA_WIDTH(24)) constant182(
    .ctrl_valid (fork22_outs_18_valid),
    .ctrl_ready (fork22_outs_18_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant182_outs),
    .outs_valid (constant182_outs_valid),
    .outs_ready (constant182_outs_ready)
  );

  handshake_constant_6 #(.DATA_WIDTH(21)) constant183(
    .ctrl_valid (fork22_outs_17_valid),
    .ctrl_ready (fork22_outs_17_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant183_outs),
    .outs_valid (constant183_outs_valid),
    .outs_ready (constant183_outs_ready)
  );

  handshake_constant_5 #(.DATA_WIDTH(18)) constant184(
    .ctrl_valid (fork22_outs_16_valid),
    .ctrl_ready (fork22_outs_16_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant184_outs),
    .outs_valid (constant184_outs_valid),
    .outs_ready (constant184_outs_ready)
  );

  handshake_constant_4 #(.DATA_WIDTH(14)) constant185(
    .ctrl_valid (fork22_outs_15_valid),
    .ctrl_ready (fork22_outs_15_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant185_outs),
    .outs_valid (constant185_outs_valid),
    .outs_ready (constant185_outs_ready)
  );

  handshake_constant_3 #(.DATA_WIDTH(12)) constant186(
    .ctrl_valid (fork22_outs_14_valid),
    .ctrl_ready (fork22_outs_14_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant186_outs),
    .outs_valid (constant186_outs_valid),
    .outs_ready (constant186_outs_ready)
  );

  handshake_constant_2 #(.DATA_WIDTH(7)) constant254(
    .ctrl_valid (fork22_outs_4_valid),
    .ctrl_ready (fork22_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant254_outs),
    .outs_valid (constant254_outs_valid),
    .outs_ready (constant254_outs_ready)
  );

  handshake_constant_1 #(.DATA_WIDTH(8)) constant188(
    .ctrl_valid (fork22_outs_13_valid),
    .ctrl_ready (fork22_outs_13_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant188_outs),
    .outs_valid (constant188_outs_valid),
    .outs_ready (constant188_outs_ready)
  );

  handshake_constant_80 #(.DATA_WIDTH(36)) constant189(
    .ctrl_valid (fork22_outs_12_valid),
    .ctrl_ready (fork22_outs_12_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant189_outs),
    .outs_valid (constant189_outs_valid),
    .outs_ready (constant189_outs_ready)
  );

  handshake_constant_81 #(.DATA_WIDTH(28)) constant255(
    .ctrl_valid (fork22_outs_3_valid),
    .ctrl_ready (fork22_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant255_outs),
    .outs_valid (constant255_outs_valid),
    .outs_ready (constant255_outs_ready)
  );

  handshake_constant_82 #(.DATA_WIDTH(30)) constant191(
    .ctrl_valid (fork22_outs_11_valid),
    .ctrl_ready (fork22_outs_11_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant191_outs),
    .outs_valid (constant191_outs_valid),
    .outs_ready (constant191_outs_ready)
  );

  handshake_constant_83 #(.DATA_WIDTH(22)) constant256(
    .ctrl_valid (fork22_outs_2_valid),
    .ctrl_ready (fork22_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant256_outs),
    .outs_valid (constant256_outs_valid),
    .outs_ready (constant256_outs_ready)
  );

  handshake_constant_84 #(.DATA_WIDTH(24)) constant193(
    .ctrl_valid (fork22_outs_10_valid),
    .ctrl_ready (fork22_outs_10_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant193_outs),
    .outs_valid (constant193_outs_valid),
    .outs_ready (constant193_outs_ready)
  );

  handshake_constant_85 #(.DATA_WIDTH(15)) constant257(
    .ctrl_valid (fork22_outs_1_valid),
    .ctrl_ready (fork22_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant257_outs),
    .outs_valid (constant257_outs_valid),
    .outs_ready (constant257_outs_ready)
  );

  handshake_constant_86 #(.DATA_WIDTH(18)) constant195(
    .ctrl_valid (fork22_outs_9_valid),
    .ctrl_ready (fork22_outs_9_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant195_outs),
    .outs_valid (constant195_outs_valid),
    .outs_ready (constant195_outs_ready)
  );

  handshake_constant_87 #(.DATA_WIDTH(8)) constant258(
    .ctrl_valid (fork22_outs_0_valid),
    .ctrl_ready (fork22_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant258_outs),
    .outs_valid (constant258_outs_valid),
    .outs_ready (constant258_outs_ready)
  );

  handshake_constant_88 #(.DATA_WIDTH(12)) constant197(
    .ctrl_valid (fork22_outs_8_valid),
    .ctrl_ready (fork22_outs_8_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant197_outs),
    .outs_valid (constant197_outs_valid),
    .outs_ready (constant197_outs_ready)
  );

  handshake_constant_89 #(.DATA_WIDTH(8)) constant198(
    .ctrl_valid (fork22_outs_7_valid),
    .ctrl_ready (fork22_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant198_outs),
    .outs_valid (constant198_outs_valid),
    .outs_ready (constant198_outs_ready)
  );

  handshake_constant_90 #(.DATA_WIDTH(8)) constant199(
    .ctrl_valid (fork22_outs_6_valid),
    .ctrl_ready (fork22_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant199_outs),
    .outs_valid (constant199_outs_valid),
    .outs_ready (constant199_outs_ready)
  );

  source source8(
    .clk (clk),
    .rst (rst),
    .outs_valid (source8_outs_valid),
    .outs_ready (source8_outs_ready)
  );

  handshake_constant_91 #(.DATA_WIDTH(4)) constant259(
    .ctrl_valid (source8_outs_valid),
    .ctrl_ready (source8_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant259_outs),
    .outs_valid (constant259_outs_valid),
    .outs_ready (constant259_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(4)) cmpi7(
    .lhs (extsi137_outs),
    .lhs_valid (extsi137_outs_valid),
    .lhs_ready (extsi137_outs_ready),
    .rhs (constant259_outs),
    .rhs_valid (constant259_outs_valid),
    .rhs_ready (constant259_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi7_result),
    .result_valid (cmpi7_result_valid),
    .result_ready (cmpi7_result_ready)
  );

  fork_type #(.SIZE(24), .DATA_TYPE(1)) fork23(
    .ins (cmpi7_result),
    .ins_valid (cmpi7_result_valid),
    .ins_ready (cmpi7_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork23_outs_23, fork23_outs_22, fork23_outs_21, fork23_outs_20, fork23_outs_19, fork23_outs_18, fork23_outs_17, fork23_outs_16, fork23_outs_15, fork23_outs_14, fork23_outs_13, fork23_outs_12, fork23_outs_11, fork23_outs_10, fork23_outs_9, fork23_outs_8, fork23_outs_7, fork23_outs_6, fork23_outs_5, fork23_outs_4, fork23_outs_3, fork23_outs_2, fork23_outs_1, fork23_outs_0}),
    .outs_valid ({fork23_outs_23_valid, fork23_outs_22_valid, fork23_outs_21_valid, fork23_outs_20_valid, fork23_outs_19_valid, fork23_outs_18_valid, fork23_outs_17_valid, fork23_outs_16_valid, fork23_outs_15_valid, fork23_outs_14_valid, fork23_outs_13_valid, fork23_outs_12_valid, fork23_outs_11_valid, fork23_outs_10_valid, fork23_outs_9_valid, fork23_outs_8_valid, fork23_outs_7_valid, fork23_outs_6_valid, fork23_outs_5_valid, fork23_outs_4_valid, fork23_outs_3_valid, fork23_outs_2_valid, fork23_outs_1_valid, fork23_outs_0_valid}),
    .outs_ready ({fork23_outs_23_ready, fork23_outs_22_ready, fork23_outs_21_ready, fork23_outs_20_ready, fork23_outs_19_ready, fork23_outs_18_ready, fork23_outs_17_ready, fork23_outs_16_ready, fork23_outs_15_ready, fork23_outs_14_ready, fork23_outs_13_ready, fork23_outs_12_ready, fork23_outs_11_ready, fork23_outs_10_ready, fork23_outs_9_ready, fork23_outs_8_ready, fork23_outs_7_ready, fork23_outs_6_ready, fork23_outs_5_ready, fork23_outs_4_ready, fork23_outs_3_ready, fork23_outs_2_ready, fork23_outs_1_ready, fork23_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(36)) cond_br106(
    .condition (fork23_outs_17),
    .condition_valid (fork23_outs_17_valid),
    .condition_ready (fork23_outs_17_ready),
    .data (constant189_outs),
    .data_valid (constant189_outs_valid),
    .data_ready (constant189_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br106_trueOut),
    .trueOut_valid (cond_br106_trueOut_valid),
    .trueOut_ready (cond_br106_trueOut_ready),
    .falseOut (cond_br106_falseOut),
    .falseOut_valid (cond_br106_falseOut_valid),
    .falseOut_ready (cond_br106_falseOut_ready)
  );

  sink #(.DATA_TYPE(36)) sink91(
    .ins (cond_br106_falseOut),
    .ins_valid (cond_br106_falseOut_valid),
    .ins_ready (cond_br106_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(28)) cond_br107(
    .condition (fork23_outs_23),
    .condition_valid (fork23_outs_23_valid),
    .condition_ready (fork23_outs_23_ready),
    .data (constant255_outs),
    .data_valid (constant255_outs_valid),
    .data_ready (constant255_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br107_trueOut),
    .trueOut_valid (cond_br107_trueOut_valid),
    .trueOut_ready (cond_br107_trueOut_ready),
    .falseOut (cond_br107_falseOut),
    .falseOut_valid (cond_br107_falseOut_valid),
    .falseOut_ready (cond_br107_falseOut_ready)
  );

  sink #(.DATA_TYPE(28)) sink92(
    .ins (cond_br107_falseOut),
    .ins_valid (cond_br107_falseOut_valid),
    .ins_ready (cond_br107_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(28), .OUTPUT_TYPE(34)) extsi138(
    .ins (cond_br107_trueOut),
    .ins_valid (cond_br107_trueOut_valid),
    .ins_ready (cond_br107_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi138_outs),
    .outs_valid (extsi138_outs_valid),
    .outs_ready (extsi138_outs_ready)
  );

  cond_br #(.DATA_TYPE(30)) cond_br108(
    .condition (fork23_outs_16),
    .condition_valid (fork23_outs_16_valid),
    .condition_ready (fork23_outs_16_ready),
    .data (constant191_outs),
    .data_valid (constant191_outs_valid),
    .data_ready (constant191_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br108_trueOut),
    .trueOut_valid (cond_br108_trueOut_valid),
    .trueOut_ready (cond_br108_trueOut_ready),
    .falseOut (cond_br108_falseOut),
    .falseOut_valid (cond_br108_falseOut_valid),
    .falseOut_ready (cond_br108_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink93(
    .ins (cond_br108_falseOut),
    .ins_valid (cond_br108_falseOut_valid),
    .ins_ready (cond_br108_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(22)) cond_br109(
    .condition (fork23_outs_22),
    .condition_valid (fork23_outs_22_valid),
    .condition_ready (fork23_outs_22_ready),
    .data (constant256_outs),
    .data_valid (constant256_outs_valid),
    .data_ready (constant256_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br109_trueOut),
    .trueOut_valid (cond_br109_trueOut_valid),
    .trueOut_ready (cond_br109_trueOut_ready),
    .falseOut (cond_br109_falseOut),
    .falseOut_valid (cond_br109_falseOut_valid),
    .falseOut_ready (cond_br109_falseOut_ready)
  );

  sink #(.DATA_TYPE(22)) sink94(
    .ins (cond_br109_falseOut),
    .ins_valid (cond_br109_falseOut_valid),
    .ins_ready (cond_br109_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(22), .OUTPUT_TYPE(27)) extsi139(
    .ins (cond_br109_trueOut),
    .ins_valid (cond_br109_trueOut_valid),
    .ins_ready (cond_br109_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi139_outs),
    .outs_valid (extsi139_outs_valid),
    .outs_ready (extsi139_outs_ready)
  );

  cond_br #(.DATA_TYPE(24)) cond_br110(
    .condition (fork23_outs_15),
    .condition_valid (fork23_outs_15_valid),
    .condition_ready (fork23_outs_15_ready),
    .data (constant193_outs),
    .data_valid (constant193_outs_valid),
    .data_ready (constant193_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br110_trueOut),
    .trueOut_valid (cond_br110_trueOut_valid),
    .trueOut_ready (cond_br110_trueOut_ready),
    .falseOut (cond_br110_falseOut),
    .falseOut_valid (cond_br110_falseOut_valid),
    .falseOut_ready (cond_br110_falseOut_ready)
  );

  sink #(.DATA_TYPE(24)) sink95(
    .ins (cond_br110_falseOut),
    .ins_valid (cond_br110_falseOut_valid),
    .ins_ready (cond_br110_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(15)) cond_br111(
    .condition (fork23_outs_21),
    .condition_valid (fork23_outs_21_valid),
    .condition_ready (fork23_outs_21_ready),
    .data (constant257_outs),
    .data_valid (constant257_outs_valid),
    .data_ready (constant257_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br111_trueOut),
    .trueOut_valid (cond_br111_trueOut_valid),
    .trueOut_ready (cond_br111_trueOut_ready),
    .falseOut (cond_br111_falseOut),
    .falseOut_valid (cond_br111_falseOut_valid),
    .falseOut_ready (cond_br111_falseOut_ready)
  );

  sink #(.DATA_TYPE(15)) sink96(
    .ins (cond_br111_falseOut),
    .ins_valid (cond_br111_falseOut_valid),
    .ins_ready (cond_br111_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(15), .OUTPUT_TYPE(21)) extsi140(
    .ins (cond_br111_trueOut),
    .ins_valid (cond_br111_trueOut_valid),
    .ins_ready (cond_br111_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi140_outs),
    .outs_valid (extsi140_outs_valid),
    .outs_ready (extsi140_outs_ready)
  );

  cond_br #(.DATA_TYPE(18)) cond_br112(
    .condition (fork23_outs_14),
    .condition_valid (fork23_outs_14_valid),
    .condition_ready (fork23_outs_14_ready),
    .data (constant195_outs),
    .data_valid (constant195_outs_valid),
    .data_ready (constant195_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br112_trueOut),
    .trueOut_valid (cond_br112_trueOut_valid),
    .trueOut_ready (cond_br112_trueOut_ready),
    .falseOut (cond_br112_falseOut),
    .falseOut_valid (cond_br112_falseOut_valid),
    .falseOut_ready (cond_br112_falseOut_ready)
  );

  sink #(.DATA_TYPE(18)) sink97(
    .ins (cond_br112_falseOut),
    .ins_valid (cond_br112_falseOut_valid),
    .ins_ready (cond_br112_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(8)) cond_br113(
    .condition (fork23_outs_20),
    .condition_valid (fork23_outs_20_valid),
    .condition_ready (fork23_outs_20_ready),
    .data (constant258_outs),
    .data_valid (constant258_outs_valid),
    .data_ready (constant258_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br113_trueOut),
    .trueOut_valid (cond_br113_trueOut_valid),
    .trueOut_ready (cond_br113_trueOut_ready),
    .falseOut (cond_br113_falseOut),
    .falseOut_valid (cond_br113_falseOut_valid),
    .falseOut_ready (cond_br113_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink98(
    .ins (cond_br113_falseOut),
    .ins_valid (cond_br113_falseOut_valid),
    .ins_ready (cond_br113_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(14)) extsi141(
    .ins (cond_br113_trueOut),
    .ins_valid (cond_br113_trueOut_valid),
    .ins_ready (cond_br113_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi141_outs),
    .outs_valid (extsi141_outs_valid),
    .outs_ready (extsi141_outs_ready)
  );

  cond_br #(.DATA_TYPE(12)) cond_br114(
    .condition (fork23_outs_13),
    .condition_valid (fork23_outs_13_valid),
    .condition_ready (fork23_outs_13_ready),
    .data (constant197_outs),
    .data_valid (constant197_outs_valid),
    .data_ready (constant197_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br114_trueOut),
    .trueOut_valid (cond_br114_trueOut_valid),
    .trueOut_ready (cond_br114_trueOut_ready),
    .falseOut (cond_br114_falseOut),
    .falseOut_valid (cond_br114_falseOut_valid),
    .falseOut_ready (cond_br114_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink99(
    .ins (cond_br114_falseOut),
    .ins_valid (cond_br114_falseOut_valid),
    .ins_ready (cond_br114_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(8)) cond_br115(
    .condition (fork23_outs_12),
    .condition_valid (fork23_outs_12_valid),
    .condition_ready (fork23_outs_12_ready),
    .data (constant198_outs),
    .data_valid (constant198_outs_valid),
    .data_ready (constant198_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br115_trueOut),
    .trueOut_valid (cond_br115_trueOut_valid),
    .trueOut_ready (cond_br115_trueOut_ready),
    .falseOut (cond_br115_falseOut),
    .falseOut_valid (cond_br115_falseOut_valid),
    .falseOut_ready (cond_br115_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink100(
    .ins (cond_br115_falseOut),
    .ins_valid (cond_br115_falseOut_valid),
    .ins_ready (cond_br115_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(8)) cond_br116(
    .condition (fork23_outs_11),
    .condition_valid (fork23_outs_11_valid),
    .condition_ready (fork23_outs_11_ready),
    .data (constant199_outs),
    .data_valid (constant199_outs_valid),
    .data_ready (constant199_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br116_trueOut),
    .trueOut_valid (cond_br116_trueOut_valid),
    .trueOut_ready (cond_br116_trueOut_ready),
    .falseOut (cond_br116_falseOut),
    .falseOut_valid (cond_br116_falseOut_valid),
    .falseOut_ready (cond_br116_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink101(
    .ins (cond_br116_falseOut),
    .ins_valid (cond_br116_falseOut_valid),
    .ins_ready (cond_br116_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer36(
    .ins (cond_br103_falseOut),
    .ins_valid (cond_br103_falseOut_valid),
    .ins_ready (cond_br103_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer36_outs),
    .outs_valid (buffer36_outs_valid),
    .outs_ready (buffer36_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer37(
    .ins (buffer36_outs),
    .ins_valid (buffer36_outs_valid),
    .ins_ready (buffer36_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer37_outs),
    .outs_valid (buffer37_outs_valid),
    .outs_ready (buffer37_outs_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br117(
    .condition (fork23_outs_0),
    .condition_valid (fork23_outs_0_valid),
    .condition_ready (fork23_outs_0_ready),
    .data (buffer37_outs),
    .data_valid (buffer37_outs_valid),
    .data_ready (buffer37_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br117_trueOut),
    .trueOut_valid (cond_br117_trueOut_valid),
    .trueOut_ready (cond_br117_trueOut_ready),
    .falseOut (cond_br117_falseOut),
    .falseOut_valid (cond_br117_falseOut_valid),
    .falseOut_ready (cond_br117_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink102(
    .ins (cond_br117_falseOut),
    .ins_valid (cond_br117_falseOut_valid),
    .ins_ready (cond_br117_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork24(
    .ins (cond_br117_trueOut),
    .ins_valid (cond_br117_trueOut_valid),
    .ins_ready (cond_br117_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork24_outs_1, fork24_outs_0}),
    .outs_valid ({fork24_outs_1_valid, fork24_outs_0_valid}),
    .outs_ready ({fork24_outs_1_ready, fork24_outs_0_ready})
  );

  cond_br_dataless cond_br118(
    .condition (fork23_outs_10),
    .condition_valid (fork23_outs_10_valid),
    .condition_ready (fork23_outs_10_ready),
    .data_valid (fork22_outs_22_valid),
    .data_ready (fork22_outs_22_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br118_trueOut_valid),
    .trueOut_ready (cond_br118_trueOut_ready),
    .falseOut_valid (cond_br118_falseOut_valid),
    .falseOut_ready (cond_br118_falseOut_ready)
  );

  sink_dataless sink103(
    .ins_valid (cond_br118_falseOut_valid),
    .ins_ready (cond_br118_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  fork_dataless #(.SIZE(2)) fork25(
    .ins_valid (cond_br118_trueOut_valid),
    .ins_ready (cond_br118_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork25_outs_1_valid, fork25_outs_0_valid}),
    .outs_ready ({fork25_outs_1_ready, fork25_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(34)) cond_br119(
    .condition (fork23_outs_19),
    .condition_valid (fork23_outs_19_valid),
    .condition_ready (fork23_outs_19_ready),
    .data (constant253_outs),
    .data_valid (constant253_outs_valid),
    .data_ready (constant253_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br119_trueOut),
    .trueOut_valid (cond_br119_trueOut_valid),
    .trueOut_ready (cond_br119_trueOut_ready),
    .falseOut (cond_br119_falseOut),
    .falseOut_valid (cond_br119_falseOut_valid),
    .falseOut_ready (cond_br119_falseOut_ready)
  );

  sink #(.DATA_TYPE(34)) sink104(
    .ins (cond_br119_falseOut),
    .ins_valid (cond_br119_falseOut_valid),
    .ins_ready (cond_br119_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(34), .OUTPUT_TYPE(36)) extsi142(
    .ins (cond_br119_trueOut),
    .ins_valid (cond_br119_trueOut_valid),
    .ins_ready (cond_br119_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi142_outs),
    .outs_valid (extsi142_outs_valid),
    .outs_ready (extsi142_outs_ready)
  );

  cond_br #(.DATA_TYPE(34)) cond_br120(
    .condition (fork23_outs_9),
    .condition_valid (fork23_outs_9_valid),
    .condition_ready (fork23_outs_9_ready),
    .data (constant179_outs),
    .data_valid (constant179_outs_valid),
    .data_ready (constant179_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br120_trueOut),
    .trueOut_valid (cond_br120_trueOut_valid),
    .trueOut_ready (cond_br120_trueOut_ready),
    .falseOut (cond_br120_falseOut),
    .falseOut_valid (cond_br120_falseOut_valid),
    .falseOut_ready (cond_br120_falseOut_ready)
  );

  sink #(.DATA_TYPE(34)) sink105(
    .ins (cond_br120_falseOut),
    .ins_valid (cond_br120_falseOut_valid),
    .ins_ready (cond_br120_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(30)) cond_br121(
    .condition (fork23_outs_8),
    .condition_valid (fork23_outs_8_valid),
    .condition_ready (fork23_outs_8_ready),
    .data (constant180_outs),
    .data_valid (constant180_outs_valid),
    .data_ready (constant180_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br121_trueOut),
    .trueOut_valid (cond_br121_trueOut_valid),
    .trueOut_ready (cond_br121_trueOut_ready),
    .falseOut (cond_br121_falseOut),
    .falseOut_valid (cond_br121_falseOut_valid),
    .falseOut_ready (cond_br121_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink106(
    .ins (cond_br121_falseOut),
    .ins_valid (cond_br121_falseOut_valid),
    .ins_ready (cond_br121_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br122(
    .condition (fork23_outs_7),
    .condition_valid (fork23_outs_7_valid),
    .condition_ready (fork23_outs_7_ready),
    .data (constant181_outs),
    .data_valid (constant181_outs_valid),
    .data_ready (constant181_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br122_trueOut),
    .trueOut_valid (cond_br122_trueOut_valid),
    .trueOut_ready (cond_br122_trueOut_ready),
    .falseOut (cond_br122_falseOut),
    .falseOut_valid (cond_br122_falseOut_valid),
    .falseOut_ready (cond_br122_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink107(
    .ins (cond_br122_falseOut),
    .ins_valid (cond_br122_falseOut_valid),
    .ins_ready (cond_br122_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(24)) cond_br123(
    .condition (fork23_outs_6),
    .condition_valid (fork23_outs_6_valid),
    .condition_ready (fork23_outs_6_ready),
    .data (constant182_outs),
    .data_valid (constant182_outs_valid),
    .data_ready (constant182_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br123_trueOut),
    .trueOut_valid (cond_br123_trueOut_valid),
    .trueOut_ready (cond_br123_trueOut_ready),
    .falseOut (cond_br123_falseOut),
    .falseOut_valid (cond_br123_falseOut_valid),
    .falseOut_ready (cond_br123_falseOut_ready)
  );

  sink #(.DATA_TYPE(24)) sink108(
    .ins (cond_br123_falseOut),
    .ins_valid (cond_br123_falseOut_valid),
    .ins_ready (cond_br123_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(21)) cond_br124(
    .condition (fork23_outs_5),
    .condition_valid (fork23_outs_5_valid),
    .condition_ready (fork23_outs_5_ready),
    .data (constant183_outs),
    .data_valid (constant183_outs_valid),
    .data_ready (constant183_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br124_trueOut),
    .trueOut_valid (cond_br124_trueOut_valid),
    .trueOut_ready (cond_br124_trueOut_ready),
    .falseOut (cond_br124_falseOut),
    .falseOut_valid (cond_br124_falseOut_valid),
    .falseOut_ready (cond_br124_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink109(
    .ins (cond_br124_falseOut),
    .ins_valid (cond_br124_falseOut_valid),
    .ins_ready (cond_br124_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(18)) cond_br125(
    .condition (fork23_outs_4),
    .condition_valid (fork23_outs_4_valid),
    .condition_ready (fork23_outs_4_ready),
    .data (constant184_outs),
    .data_valid (constant184_outs_valid),
    .data_ready (constant184_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br125_trueOut),
    .trueOut_valid (cond_br125_trueOut_valid),
    .trueOut_ready (cond_br125_trueOut_ready),
    .falseOut (cond_br125_falseOut),
    .falseOut_valid (cond_br125_falseOut_valid),
    .falseOut_ready (cond_br125_falseOut_ready)
  );

  sink #(.DATA_TYPE(18)) sink110(
    .ins (cond_br125_falseOut),
    .ins_valid (cond_br125_falseOut_valid),
    .ins_ready (cond_br125_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(14)) cond_br126(
    .condition (fork23_outs_3),
    .condition_valid (fork23_outs_3_valid),
    .condition_ready (fork23_outs_3_ready),
    .data (constant185_outs),
    .data_valid (constant185_outs_valid),
    .data_ready (constant185_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br126_trueOut),
    .trueOut_valid (cond_br126_trueOut_valid),
    .trueOut_ready (cond_br126_trueOut_ready),
    .falseOut (cond_br126_falseOut),
    .falseOut_valid (cond_br126_falseOut_valid),
    .falseOut_ready (cond_br126_falseOut_ready)
  );

  sink #(.DATA_TYPE(14)) sink111(
    .ins (cond_br126_falseOut),
    .ins_valid (cond_br126_falseOut_valid),
    .ins_ready (cond_br126_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br127(
    .condition (fork23_outs_2),
    .condition_valid (fork23_outs_2_valid),
    .condition_ready (fork23_outs_2_ready),
    .data (constant186_outs),
    .data_valid (constant186_outs_valid),
    .data_ready (constant186_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br127_trueOut),
    .trueOut_valid (cond_br127_trueOut_valid),
    .trueOut_ready (cond_br127_trueOut_ready),
    .falseOut (cond_br127_falseOut),
    .falseOut_valid (cond_br127_falseOut_valid),
    .falseOut_ready (cond_br127_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink112(
    .ins (cond_br127_falseOut),
    .ins_valid (cond_br127_falseOut_valid),
    .ins_ready (cond_br127_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br128(
    .condition (fork23_outs_18),
    .condition_valid (fork23_outs_18_valid),
    .condition_ready (fork23_outs_18_ready),
    .data (constant254_outs),
    .data_valid (constant254_outs_valid),
    .data_ready (constant254_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br128_trueOut),
    .trueOut_valid (cond_br128_trueOut_valid),
    .trueOut_ready (cond_br128_trueOut_ready),
    .falseOut (cond_br128_falseOut),
    .falseOut_valid (cond_br128_falseOut_valid),
    .falseOut_ready (cond_br128_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink113(
    .ins (cond_br128_falseOut),
    .ins_valid (cond_br128_falseOut_valid),
    .ins_ready (cond_br128_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(8)) extsi143(
    .ins (cond_br128_trueOut),
    .ins_valid (cond_br128_trueOut_valid),
    .ins_ready (cond_br128_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi143_outs),
    .outs_valid (extsi143_outs_valid),
    .outs_ready (extsi143_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br129(
    .condition (fork23_outs_1),
    .condition_valid (fork23_outs_1_valid),
    .condition_ready (fork23_outs_1_ready),
    .data (constant188_outs),
    .data_valid (constant188_outs_valid),
    .data_ready (constant188_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br129_trueOut),
    .trueOut_valid (cond_br129_trueOut_valid),
    .trueOut_ready (cond_br129_trueOut_ready),
    .falseOut (cond_br129_falseOut),
    .falseOut_valid (cond_br129_falseOut_valid),
    .falseOut_ready (cond_br129_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink114(
    .ins (cond_br129_falseOut),
    .ins_valid (cond_br129_falseOut_valid),
    .ins_ready (cond_br129_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  mux #(.SIZE(9), .DATA_TYPE(36), .SELECT_TYPE(4)) mux0(
    .index (fork27_outs_11),
    .index_valid (fork27_outs_11_valid),
    .index_ready (fork27_outs_11_ready),
    .ins ({extsi142_outs, cond_br106_trueOut, cond_br92_trueOut, cond_br78_trueOut, cond_br64_trueOut, cond_br50_trueOut, cond_br36_trueOut, extsi103_outs, extsi100_outs}),
    .ins_valid ({extsi142_outs_valid, cond_br106_trueOut_valid, cond_br92_trueOut_valid, cond_br78_trueOut_valid, cond_br64_trueOut_valid, cond_br50_trueOut_valid, cond_br36_trueOut_valid, extsi103_outs_valid, extsi100_outs_valid}),
    .ins_ready ({extsi142_outs_ready, cond_br106_trueOut_ready, cond_br92_trueOut_ready, cond_br78_trueOut_ready, cond_br64_trueOut_ready, cond_br50_trueOut_ready, cond_br36_trueOut_ready, extsi103_outs_ready, extsi100_outs_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux0_outs),
    .outs_valid (mux0_outs_valid),
    .outs_ready (mux0_outs_ready)
  );

  mux #(.SIZE(9), .DATA_TYPE(34), .SELECT_TYPE(4)) mux1(
    .index (fork27_outs_10),
    .index_valid (fork27_outs_10_valid),
    .index_ready (fork27_outs_10_ready),
    .ins ({cond_br120_trueOut, extsi138_outs, extsi132_outs, extsi126_outs, extsi119_outs, extsi113_outs, extsi106_outs, extsi104_outs, cond_br9_trueOut}),
    .ins_valid ({cond_br120_trueOut_valid, extsi138_outs_valid, extsi132_outs_valid, extsi126_outs_valid, extsi119_outs_valid, extsi113_outs_valid, extsi106_outs_valid, extsi104_outs_valid, cond_br9_trueOut_valid}),
    .ins_ready ({cond_br120_trueOut_ready, extsi138_outs_ready, extsi132_outs_ready, extsi126_outs_ready, extsi119_outs_ready, extsi113_outs_ready, extsi106_outs_ready, extsi104_outs_ready, cond_br9_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux1_outs),
    .outs_valid (mux1_outs_valid),
    .outs_ready (mux1_outs_ready)
  );

  mux #(.SIZE(9), .DATA_TYPE(30), .SELECT_TYPE(4)) mux2(
    .index (fork27_outs_9),
    .index_valid (fork27_outs_9_valid),
    .index_ready (fork27_outs_9_ready),
    .ins ({cond_br121_trueOut, cond_br108_trueOut, cond_br94_trueOut, cond_br80_trueOut, cond_br66_trueOut, cond_br52_trueOut, cond_br38_trueOut, cond_br24_trueOut, cond_br10_trueOut}),
    .ins_valid ({cond_br121_trueOut_valid, cond_br108_trueOut_valid, cond_br94_trueOut_valid, cond_br80_trueOut_valid, cond_br66_trueOut_valid, cond_br52_trueOut_valid, cond_br38_trueOut_valid, cond_br24_trueOut_valid, cond_br10_trueOut_valid}),
    .ins_ready ({cond_br121_trueOut_ready, cond_br108_trueOut_ready, cond_br94_trueOut_ready, cond_br80_trueOut_ready, cond_br66_trueOut_ready, cond_br52_trueOut_ready, cond_br38_trueOut_ready, cond_br24_trueOut_ready, cond_br10_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux2_outs),
    .outs_valid (mux2_outs_valid),
    .outs_ready (mux2_outs_ready)
  );

  mux #(.SIZE(9), .DATA_TYPE(27), .SELECT_TYPE(4)) mux3(
    .index (fork27_outs_8),
    .index_valid (fork27_outs_8_valid),
    .index_ready (fork27_outs_8_ready),
    .ins ({cond_br122_trueOut, extsi139_outs, extsi133_outs, extsi127_outs, extsi120_outs, extsi114_outs, extsi107_outs, cond_br25_trueOut, cond_br11_trueOut}),
    .ins_valid ({cond_br122_trueOut_valid, extsi139_outs_valid, extsi133_outs_valid, extsi127_outs_valid, extsi120_outs_valid, extsi114_outs_valid, extsi107_outs_valid, cond_br25_trueOut_valid, cond_br11_trueOut_valid}),
    .ins_ready ({cond_br122_trueOut_ready, extsi139_outs_ready, extsi133_outs_ready, extsi127_outs_ready, extsi120_outs_ready, extsi114_outs_ready, extsi107_outs_ready, cond_br25_trueOut_ready, cond_br11_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux3_outs),
    .outs_valid (mux3_outs_valid),
    .outs_ready (mux3_outs_ready)
  );

  mux #(.SIZE(9), .DATA_TYPE(24), .SELECT_TYPE(4)) mux4(
    .index (fork27_outs_7),
    .index_valid (fork27_outs_7_valid),
    .index_ready (fork27_outs_7_ready),
    .ins ({cond_br123_trueOut, cond_br110_trueOut, cond_br96_trueOut, cond_br82_trueOut, cond_br68_trueOut, cond_br54_trueOut, extsi108_outs, cond_br26_trueOut, cond_br12_trueOut}),
    .ins_valid ({cond_br123_trueOut_valid, cond_br110_trueOut_valid, cond_br96_trueOut_valid, cond_br82_trueOut_valid, cond_br68_trueOut_valid, cond_br54_trueOut_valid, extsi108_outs_valid, cond_br26_trueOut_valid, cond_br12_trueOut_valid}),
    .ins_ready ({cond_br123_trueOut_ready, cond_br110_trueOut_ready, cond_br96_trueOut_ready, cond_br82_trueOut_ready, cond_br68_trueOut_ready, cond_br54_trueOut_ready, extsi108_outs_ready, cond_br26_trueOut_ready, cond_br12_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux4_outs),
    .outs_valid (mux4_outs_valid),
    .outs_ready (mux4_outs_ready)
  );

  mux #(.SIZE(9), .DATA_TYPE(21), .SELECT_TYPE(4)) mux5(
    .index (fork27_outs_6),
    .index_valid (fork27_outs_6_valid),
    .index_ready (fork27_outs_6_ready),
    .ins ({cond_br124_trueOut, extsi140_outs, extsi134_outs, extsi128_outs, extsi121_outs, cond_br55_trueOut, cond_br41_trueOut, cond_br27_trueOut, cond_br13_trueOut}),
    .ins_valid ({cond_br124_trueOut_valid, extsi140_outs_valid, extsi134_outs_valid, extsi128_outs_valid, extsi121_outs_valid, cond_br55_trueOut_valid, cond_br41_trueOut_valid, cond_br27_trueOut_valid, cond_br13_trueOut_valid}),
    .ins_ready ({cond_br124_trueOut_ready, extsi140_outs_ready, extsi134_outs_ready, extsi128_outs_ready, extsi121_outs_ready, cond_br55_trueOut_ready, cond_br41_trueOut_ready, cond_br27_trueOut_ready, cond_br13_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux5_outs),
    .outs_valid (mux5_outs_valid),
    .outs_ready (mux5_outs_ready)
  );

  mux #(.SIZE(9), .DATA_TYPE(18), .SELECT_TYPE(4)) mux6(
    .index (fork27_outs_5),
    .index_valid (fork27_outs_5_valid),
    .index_ready (fork27_outs_5_ready),
    .ins ({cond_br125_trueOut, cond_br112_trueOut, cond_br98_trueOut, cond_br84_trueOut, extsi122_outs, extsi115_outs, extsi109_outs, cond_br28_trueOut, cond_br14_trueOut}),
    .ins_valid ({cond_br125_trueOut_valid, cond_br112_trueOut_valid, cond_br98_trueOut_valid, cond_br84_trueOut_valid, extsi122_outs_valid, extsi115_outs_valid, extsi109_outs_valid, cond_br28_trueOut_valid, cond_br14_trueOut_valid}),
    .ins_ready ({cond_br125_trueOut_ready, cond_br112_trueOut_ready, cond_br98_trueOut_ready, cond_br84_trueOut_ready, extsi122_outs_ready, extsi115_outs_ready, extsi109_outs_ready, cond_br28_trueOut_ready, cond_br14_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux6_outs),
    .outs_valid (mux6_outs_valid),
    .outs_ready (mux6_outs_ready)
  );

  mux #(.SIZE(9), .DATA_TYPE(14), .SELECT_TYPE(4)) mux7(
    .index (fork27_outs_4),
    .index_valid (fork27_outs_4_valid),
    .index_ready (fork27_outs_4_ready),
    .ins ({cond_br126_trueOut, extsi141_outs, extsi135_outs, cond_br85_trueOut, cond_br71_trueOut, cond_br57_trueOut, extsi110_outs, cond_br29_trueOut, cond_br15_trueOut}),
    .ins_valid ({cond_br126_trueOut_valid, extsi141_outs_valid, extsi135_outs_valid, cond_br85_trueOut_valid, cond_br71_trueOut_valid, cond_br57_trueOut_valid, extsi110_outs_valid, cond_br29_trueOut_valid, cond_br15_trueOut_valid}),
    .ins_ready ({cond_br126_trueOut_ready, extsi141_outs_ready, extsi135_outs_ready, cond_br85_trueOut_ready, cond_br71_trueOut_ready, cond_br57_trueOut_ready, extsi110_outs_ready, cond_br29_trueOut_ready, cond_br15_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux7_outs),
    .outs_valid (mux7_outs_valid),
    .outs_ready (mux7_outs_ready)
  );

  mux #(.SIZE(9), .DATA_TYPE(12), .SELECT_TYPE(4)) mux8(
    .index (fork27_outs_3),
    .index_valid (fork27_outs_3_valid),
    .index_ready (fork27_outs_3_ready),
    .ins ({cond_br127_trueOut, cond_br114_trueOut, cond_br100_trueOut, extsi129_outs, cond_br72_trueOut, cond_br58_trueOut, cond_br44_trueOut, extsi105_outs, cond_br16_trueOut}),
    .ins_valid ({cond_br127_trueOut_valid, cond_br114_trueOut_valid, cond_br100_trueOut_valid, extsi129_outs_valid, cond_br72_trueOut_valid, cond_br58_trueOut_valid, cond_br44_trueOut_valid, extsi105_outs_valid, cond_br16_trueOut_valid}),
    .ins_ready ({cond_br127_trueOut_ready, cond_br114_trueOut_ready, cond_br100_trueOut_ready, extsi129_outs_ready, cond_br72_trueOut_ready, cond_br58_trueOut_ready, cond_br44_trueOut_ready, extsi105_outs_ready, cond_br16_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux8_outs),
    .outs_valid (mux8_outs_valid),
    .outs_ready (mux8_outs_ready)
  );

  mux #(.SIZE(9), .DATA_TYPE(8), .SELECT_TYPE(4)) mux9(
    .index (fork27_outs_2),
    .index_valid (fork27_outs_2_valid),
    .index_ready (fork27_outs_2_ready),
    .ins ({extsi143_outs, cond_br115_trueOut, cond_br101_trueOut, extsi130_outs, extsi123_outs, extsi116_outs, extsi111_outs, cond_br31_trueOut, extsi101_outs}),
    .ins_valid ({extsi143_outs_valid, cond_br115_trueOut_valid, cond_br101_trueOut_valid, extsi130_outs_valid, extsi123_outs_valid, extsi116_outs_valid, extsi111_outs_valid, cond_br31_trueOut_valid, extsi101_outs_valid}),
    .ins_ready ({extsi143_outs_ready, cond_br115_trueOut_ready, cond_br101_trueOut_ready, extsi130_outs_ready, extsi123_outs_ready, extsi116_outs_ready, extsi111_outs_ready, cond_br31_trueOut_ready, extsi101_outs_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux9_outs),
    .outs_valid (mux9_outs_valid),
    .outs_ready (mux9_outs_ready)
  );

  mux #(.SIZE(9), .DATA_TYPE(8), .SELECT_TYPE(4)) mux10(
    .index (fork27_outs_1),
    .index_valid (fork27_outs_1_valid),
    .index_ready (fork27_outs_1_ready),
    .ins ({cond_br129_trueOut, cond_br116_trueOut, extsi136_outs, cond_br88_trueOut, extsi124_outs, extsi117_outs, extsi112_outs, cond_br32_trueOut, cond_br18_trueOut}),
    .ins_valid ({cond_br129_trueOut_valid, cond_br116_trueOut_valid, extsi136_outs_valid, cond_br88_trueOut_valid, extsi124_outs_valid, extsi117_outs_valid, extsi112_outs_valid, cond_br32_trueOut_valid, cond_br18_trueOut_valid}),
    .ins_ready ({cond_br129_trueOut_ready, cond_br116_trueOut_ready, extsi136_outs_ready, cond_br88_trueOut_ready, extsi124_outs_ready, extsi117_outs_ready, extsi112_outs_ready, cond_br32_trueOut_ready, cond_br18_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux10_outs),
    .outs_valid (mux10_outs_valid),
    .outs_ready (mux10_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer62(
    .ins (mux10_outs),
    .ins_valid (mux10_outs_valid),
    .ins_ready (mux10_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer62_outs),
    .outs_valid (buffer62_outs_valid),
    .outs_ready (buffer62_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer63(
    .ins (buffer62_outs),
    .ins_valid (buffer62_outs_valid),
    .ins_ready (buffer62_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer63_outs),
    .outs_valid (buffer63_outs_valid),
    .outs_ready (buffer63_outs_ready)
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(13)) extsi144(
    .ins (buffer63_outs),
    .ins_valid (buffer63_outs_valid),
    .ins_ready (buffer63_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi144_outs),
    .outs_valid (extsi144_outs_valid),
    .outs_ready (extsi144_outs_ready)
  );

  mux #(.SIZE(9), .DATA_TYPE(5), .SELECT_TYPE(4)) mux11(
    .index (fork27_outs_0),
    .index_valid (fork27_outs_0_valid),
    .index_ready (fork27_outs_0_ready),
    .ins ({fork24_outs_1, fork24_outs_0, cond_br103_trueOut, cond_br89_trueOut, cond_br75_trueOut, cond_br61_trueOut, cond_br47_trueOut, cond_br33_trueOut, cond_br19_trueOut}),
    .ins_valid ({fork24_outs_1_valid, fork24_outs_0_valid, cond_br103_trueOut_valid, cond_br89_trueOut_valid, cond_br75_trueOut_valid, cond_br61_trueOut_valid, cond_br47_trueOut_valid, cond_br33_trueOut_valid, cond_br19_trueOut_valid}),
    .ins_ready ({fork24_outs_1_ready, fork24_outs_0_ready, cond_br103_trueOut_ready, cond_br89_trueOut_ready, cond_br75_trueOut_ready, cond_br61_trueOut_ready, cond_br47_trueOut_ready, cond_br33_trueOut_ready, cond_br19_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux11_outs),
    .outs_valid (mux11_outs_valid),
    .outs_ready (mux11_outs_ready)
  );

  oehb #(.DATA_TYPE(5)) buffer64(
    .ins (mux11_outs),
    .ins_valid (mux11_outs_valid),
    .ins_ready (mux11_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer64_outs),
    .outs_valid (buffer64_outs_valid),
    .outs_ready (buffer64_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer65(
    .ins (buffer64_outs),
    .ins_valid (buffer64_outs_valid),
    .ins_ready (buffer64_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer65_outs),
    .outs_valid (buffer65_outs_valid),
    .outs_ready (buffer65_outs_ready)
  );

  fork_type #(.SIZE(10), .DATA_TYPE(5)) fork26(
    .ins (buffer65_outs),
    .ins_valid (buffer65_outs_valid),
    .ins_ready (buffer65_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork26_outs_9, fork26_outs_8, fork26_outs_7, fork26_outs_6, fork26_outs_5, fork26_outs_4, fork26_outs_3, fork26_outs_2, fork26_outs_1, fork26_outs_0}),
    .outs_valid ({fork26_outs_9_valid, fork26_outs_8_valid, fork26_outs_7_valid, fork26_outs_6_valid, fork26_outs_5_valid, fork26_outs_4_valid, fork26_outs_3_valid, fork26_outs_2_valid, fork26_outs_1_valid, fork26_outs_0_valid}),
    .outs_ready ({fork26_outs_9_ready, fork26_outs_8_ready, fork26_outs_7_ready, fork26_outs_6_ready, fork26_outs_5_ready, fork26_outs_4_ready, fork26_outs_3_ready, fork26_outs_2_ready, fork26_outs_1_ready, fork26_outs_0_ready})
  );

  control_merge_dataless #(.SIZE(9), .INDEX_TYPE(4)) control_merge7(
    .ins_valid ({fork25_outs_1_valid, fork25_outs_0_valid, cond_br104_trueOut_valid, cond_br90_trueOut_valid, cond_br76_trueOut_valid, cond_br62_trueOut_valid, cond_br48_trueOut_valid, cond_br34_trueOut_valid, cond_br20_trueOut_valid}),
    .ins_ready ({fork25_outs_1_ready, fork25_outs_0_ready, cond_br104_trueOut_ready, cond_br90_trueOut_ready, cond_br76_trueOut_ready, cond_br62_trueOut_ready, cond_br48_trueOut_ready, cond_br34_trueOut_ready, cond_br20_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs_valid (control_merge7_outs_valid),
    .outs_ready (control_merge7_outs_ready),
    .index (control_merge7_index),
    .index_valid (control_merge7_index_valid),
    .index_ready (control_merge7_index_ready)
  );

  fork_type #(.SIZE(12), .DATA_TYPE(4)) fork27(
    .ins (control_merge7_index),
    .ins_valid (control_merge7_index_valid),
    .ins_ready (control_merge7_index_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork27_outs_11, fork27_outs_10, fork27_outs_9, fork27_outs_8, fork27_outs_7, fork27_outs_6, fork27_outs_5, fork27_outs_4, fork27_outs_3, fork27_outs_2, fork27_outs_1, fork27_outs_0}),
    .outs_valid ({fork27_outs_11_valid, fork27_outs_10_valid, fork27_outs_9_valid, fork27_outs_8_valid, fork27_outs_7_valid, fork27_outs_6_valid, fork27_outs_5_valid, fork27_outs_4_valid, fork27_outs_3_valid, fork27_outs_2_valid, fork27_outs_1_valid, fork27_outs_0_valid}),
    .outs_ready ({fork27_outs_11_ready, fork27_outs_10_ready, fork27_outs_9_ready, fork27_outs_8_ready, fork27_outs_7_ready, fork27_outs_6_ready, fork27_outs_5_ready, fork27_outs_4_ready, fork27_outs_3_ready, fork27_outs_2_ready, fork27_outs_1_ready, fork27_outs_0_ready})
  );

  oehb_dataless buffer66(
    .ins_valid (control_merge7_outs_valid),
    .ins_ready (control_merge7_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer66_outs_valid),
    .outs_ready (buffer66_outs_ready)
  );

  tehb_dataless buffer67(
    .ins_valid (buffer66_outs_valid),
    .ins_ready (buffer66_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer67_outs_valid),
    .outs_ready (buffer67_outs_ready)
  );

  sink_dataless sink115(
    .ins_valid (buffer67_outs_valid),
    .ins_ready (buffer67_outs_ready),
    .clk (clk),
    .rst (rst)
  );

  source source9(
    .clk (clk),
    .rst (rst),
    .outs_valid (source9_outs_valid),
    .outs_ready (source9_outs_ready)
  );

  handshake_constant_47 #(.DATA_WIDTH(3)) constant260(
    .ctrl_valid (source9_outs_valid),
    .ctrl_ready (source9_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant260_outs),
    .outs_valid (constant260_outs_valid),
    .outs_ready (constant260_outs_ready)
  );

  fork_type #(.SIZE(10), .DATA_TYPE(3)) fork28(
    .ins (constant260_outs),
    .ins_valid (constant260_outs_valid),
    .ins_ready (constant260_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork28_outs_9, fork28_outs_8, fork28_outs_7, fork28_outs_6, fork28_outs_5, fork28_outs_4, fork28_outs_3, fork28_outs_2, fork28_outs_1, fork28_outs_0}),
    .outs_valid ({fork28_outs_9_valid, fork28_outs_8_valid, fork28_outs_7_valid, fork28_outs_6_valid, fork28_outs_5_valid, fork28_outs_4_valid, fork28_outs_3_valid, fork28_outs_2_valid, fork28_outs_1_valid, fork28_outs_0_valid}),
    .outs_ready ({fork28_outs_9_ready, fork28_outs_8_ready, fork28_outs_7_ready, fork28_outs_6_ready, fork28_outs_5_ready, fork28_outs_4_ready, fork28_outs_3_ready, fork28_outs_2_ready, fork28_outs_1_ready, fork28_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(40)) extsi88(
    .ins (fork28_outs_0),
    .ins_valid (fork28_outs_0_valid),
    .ins_ready (fork28_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi88_outs),
    .outs_valid (extsi88_outs_valid),
    .outs_ready (extsi88_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(38)) extsi89(
    .ins (fork28_outs_1),
    .ins_valid (fork28_outs_1_valid),
    .ins_ready (fork28_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi89_outs),
    .outs_valid (extsi89_outs_valid),
    .outs_ready (extsi89_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(34)) extsi90(
    .ins (fork28_outs_2),
    .ins_valid (fork28_outs_2_valid),
    .ins_ready (fork28_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi90_outs),
    .outs_valid (extsi90_outs_valid),
    .outs_ready (extsi90_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(31)) extsi91(
    .ins (fork28_outs_3),
    .ins_valid (fork28_outs_3_valid),
    .ins_ready (fork28_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi91_outs),
    .outs_valid (extsi91_outs_valid),
    .outs_ready (extsi91_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(28)) extsi92(
    .ins (fork28_outs_4),
    .ins_valid (fork28_outs_4_valid),
    .ins_ready (fork28_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi92_outs),
    .outs_valid (extsi92_outs_valid),
    .outs_ready (extsi92_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(25)) extsi93(
    .ins (fork28_outs_5),
    .ins_valid (fork28_outs_5_valid),
    .ins_ready (fork28_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi93_outs),
    .outs_valid (extsi93_outs_valid),
    .outs_ready (extsi93_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(22)) extsi94(
    .ins (fork28_outs_6),
    .ins_valid (fork28_outs_6_valid),
    .ins_ready (fork28_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi94_outs),
    .outs_valid (extsi94_outs_valid),
    .outs_ready (extsi94_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(19)) extsi95(
    .ins (fork28_outs_7),
    .ins_valid (fork28_outs_7_valid),
    .ins_ready (fork28_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi95_outs),
    .outs_valid (extsi95_outs_valid),
    .outs_ready (extsi95_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(16)) extsi96(
    .ins (fork28_outs_8),
    .ins_valid (fork28_outs_8_valid),
    .ins_ready (fork28_outs_8_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi96_outs),
    .outs_valid (extsi96_outs_valid),
    .outs_ready (extsi96_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(12)) extsi97(
    .ins (fork28_outs_9),
    .ins_valid (fork28_outs_9_valid),
    .ins_ready (fork28_outs_9_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi97_outs),
    .outs_valid (extsi97_outs_valid),
    .outs_ready (extsi97_outs_ready)
  );

  source source19(
    .clk (clk),
    .rst (rst),
    .outs_valid (source19_outs_valid),
    .outs_ready (source19_outs_ready)
  );

  handshake_constant_12 #(.DATA_WIDTH(4)) constant261(
    .ctrl_valid (source19_outs_valid),
    .ctrl_ready (source19_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant261_outs),
    .outs_valid (constant261_outs_valid),
    .outs_ready (constant261_outs_ready)
  );

  extui #(.INPUT_TYPE(4), .OUTPUT_TYPE(13)) extui0(
    .ins (constant261_outs),
    .ins_valid (constant261_outs_valid),
    .ins_ready (constant261_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extui0_outs),
    .outs_valid (extui0_outs_valid),
    .outs_ready (extui0_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(13)) extsi145(
    .ins (fork26_outs_9),
    .ins_valid (fork26_outs_9_valid),
    .ins_ready (fork26_outs_9_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi145_outs),
    .outs_valid (extsi145_outs_valid),
    .outs_ready (extsi145_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(16)) extsi146(
    .ins (fork26_outs_8),
    .ins_valid (fork26_outs_8_valid),
    .ins_ready (fork26_outs_8_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi146_outs),
    .outs_valid (extsi146_outs_valid),
    .outs_ready (extsi146_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(20)) extsi147(
    .ins (fork26_outs_7),
    .ins_valid (fork26_outs_7_valid),
    .ins_ready (fork26_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi147_outs),
    .outs_valid (extsi147_outs_valid),
    .outs_ready (extsi147_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(23)) extsi148(
    .ins (fork26_outs_6),
    .ins_valid (fork26_outs_6_valid),
    .ins_ready (fork26_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi148_outs),
    .outs_valid (extsi148_outs_valid),
    .outs_ready (extsi148_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(26)) extsi149(
    .ins (fork26_outs_5),
    .ins_valid (fork26_outs_5_valid),
    .ins_ready (fork26_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi149_outs),
    .outs_valid (extsi149_outs_valid),
    .outs_ready (extsi149_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(29)) extsi150(
    .ins (fork26_outs_4),
    .ins_valid (fork26_outs_4_valid),
    .ins_ready (fork26_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi150_outs),
    .outs_valid (extsi150_outs_valid),
    .outs_ready (extsi150_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(32)) extsi151(
    .ins (fork26_outs_3),
    .ins_valid (fork26_outs_3_valid),
    .ins_ready (fork26_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi151_outs),
    .outs_valid (extsi151_outs_valid),
    .outs_ready (extsi151_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(35)) extsi152(
    .ins (fork26_outs_2),
    .ins_valid (fork26_outs_2_valid),
    .ins_ready (fork26_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi152_outs),
    .outs_valid (extsi152_outs_valid),
    .outs_ready (extsi152_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(38)) extsi153(
    .ins (fork26_outs_1),
    .ins_valid (fork26_outs_1_valid),
    .ins_ready (fork26_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi153_outs),
    .outs_valid (extsi153_outs_valid),
    .outs_ready (extsi153_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(42)) extsi154(
    .ins (fork26_outs_0),
    .ins_valid (fork26_outs_0_valid),
    .ins_ready (fork26_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi154_outs),
    .outs_valid (extsi154_outs_valid),
    .outs_ready (extsi154_outs_ready)
  );

  muli #(.DATA_TYPE(13)) muli0(
    .lhs (extsi144_outs),
    .lhs_valid (extsi144_outs_valid),
    .lhs_ready (extsi144_outs_ready),
    .rhs (extsi145_outs),
    .rhs_valid (extsi145_outs_valid),
    .rhs_ready (extsi145_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli0_result),
    .result_valid (muli0_result_valid),
    .result_ready (muli0_result_ready)
  );

  trunci #(.INPUT_TYPE(13), .OUTPUT_TYPE(11)) trunci2(
    .ins (muli0_result),
    .ins_valid (muli0_result_valid),
    .ins_ready (muli0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci2_outs),
    .outs_valid (trunci2_outs_valid),
    .outs_ready (trunci2_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer60(
    .ins (mux9_outs),
    .ins_valid (mux9_outs_valid),
    .ins_ready (mux9_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer60_outs),
    .outs_valid (buffer60_outs_valid),
    .outs_ready (buffer60_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer61(
    .ins (buffer60_outs),
    .ins_valid (buffer60_outs_valid),
    .ins_ready (buffer60_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer61_outs),
    .outs_valid (buffer61_outs_valid),
    .outs_ready (buffer61_outs_ready)
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(12)) extsi3(
    .ins (buffer61_outs),
    .ins_valid (buffer61_outs_valid),
    .ins_ready (buffer61_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi3_outs),
    .outs_valid (extsi3_outs_valid),
    .outs_ready (extsi3_outs_ready)
  );

  shli #(.DATA_TYPE(12)) shli0(
    .lhs (extsi3_outs),
    .lhs_valid (extsi3_outs_valid),
    .lhs_ready (extsi3_outs_ready),
    .rhs (extsi97_outs),
    .rhs_valid (extsi97_outs_valid),
    .rhs_ready (extsi97_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli0_result),
    .result_valid (shli0_result_valid),
    .result_ready (shli0_result_ready)
  );

  trunci #(.INPUT_TYPE(12), .OUTPUT_TYPE(11)) trunci24(
    .ins (shli0_result),
    .ins_valid (shli0_result_valid),
    .ins_ready (shli0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci24_outs),
    .outs_valid (trunci24_outs_valid),
    .outs_ready (trunci24_outs_ready)
  );

  addi #(.DATA_TYPE(11)) addi0(
    .lhs (trunci2_outs),
    .lhs_valid (trunci2_outs_valid),
    .lhs_ready (trunci2_outs_ready),
    .rhs (trunci24_outs),
    .rhs_valid (trunci24_outs_valid),
    .rhs_ready (trunci24_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi0_result),
    .result_valid (addi0_result_valid),
    .result_ready (addi0_result_ready)
  );

  extsi #(.INPUT_TYPE(11), .OUTPUT_TYPE(16)) extsi155(
    .ins (addi0_result),
    .ins_valid (addi0_result_valid),
    .ins_ready (addi0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi155_outs),
    .outs_valid (extsi155_outs_valid),
    .outs_ready (extsi155_outs_ready)
  );

  muli #(.DATA_TYPE(16)) muli1(
    .lhs (extsi155_outs),
    .lhs_valid (extsi155_outs_valid),
    .lhs_ready (extsi155_outs_ready),
    .rhs (extsi146_outs),
    .rhs_valid (extsi146_outs_valid),
    .rhs_ready (extsi146_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli1_result),
    .result_valid (muli1_result_valid),
    .result_ready (muli1_result_ready)
  );

  trunci #(.INPUT_TYPE(16), .OUTPUT_TYPE(15)) trunci4(
    .ins (muli1_result),
    .ins_valid (muli1_result_valid),
    .ins_ready (muli1_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci4_outs),
    .outs_valid (trunci4_outs_valid),
    .outs_ready (trunci4_outs_ready)
  );

  oehb #(.DATA_TYPE(12)) buffer58(
    .ins (mux8_outs),
    .ins_valid (mux8_outs_valid),
    .ins_ready (mux8_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer58_outs),
    .outs_valid (buffer58_outs_valid),
    .outs_ready (buffer58_outs_ready)
  );

  tehb #(.DATA_TYPE(12)) buffer59(
    .ins (buffer58_outs),
    .ins_valid (buffer58_outs_valid),
    .ins_ready (buffer58_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer59_outs),
    .outs_valid (buffer59_outs_valid),
    .outs_ready (buffer59_outs_ready)
  );

  extsi #(.INPUT_TYPE(12), .OUTPUT_TYPE(16)) extsi7(
    .ins (buffer59_outs),
    .ins_valid (buffer59_outs_valid),
    .ins_ready (buffer59_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi7_outs),
    .outs_valid (extsi7_outs_valid),
    .outs_ready (extsi7_outs_ready)
  );

  shli #(.DATA_TYPE(16)) shli1(
    .lhs (extsi7_outs),
    .lhs_valid (extsi7_outs_valid),
    .lhs_ready (extsi7_outs_ready),
    .rhs (extsi96_outs),
    .rhs_valid (extsi96_outs_valid),
    .rhs_ready (extsi96_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli1_result),
    .result_valid (shli1_result_valid),
    .result_ready (shli1_result_ready)
  );

  trunci #(.INPUT_TYPE(16), .OUTPUT_TYPE(15)) trunci25(
    .ins (shli1_result),
    .ins_valid (shli1_result_valid),
    .ins_ready (shli1_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci25_outs),
    .outs_valid (trunci25_outs_valid),
    .outs_ready (trunci25_outs_ready)
  );

  addi #(.DATA_TYPE(15)) addi1(
    .lhs (trunci4_outs),
    .lhs_valid (trunci4_outs_valid),
    .lhs_ready (trunci4_outs_ready),
    .rhs (trunci25_outs),
    .rhs_valid (trunci25_outs_valid),
    .rhs_ready (trunci25_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi1_result),
    .result_valid (addi1_result_valid),
    .result_ready (addi1_result_ready)
  );

  extsi #(.INPUT_TYPE(15), .OUTPUT_TYPE(20)) extsi156(
    .ins (addi1_result),
    .ins_valid (addi1_result_valid),
    .ins_ready (addi1_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi156_outs),
    .outs_valid (extsi156_outs_valid),
    .outs_ready (extsi156_outs_ready)
  );

  muli #(.DATA_TYPE(20)) muli2(
    .lhs (extsi156_outs),
    .lhs_valid (extsi156_outs_valid),
    .lhs_ready (extsi156_outs_ready),
    .rhs (extsi147_outs),
    .rhs_valid (extsi147_outs_valid),
    .rhs_ready (extsi147_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli2_result),
    .result_valid (muli2_result_valid),
    .result_ready (muli2_result_ready)
  );

  trunci #(.INPUT_TYPE(20), .OUTPUT_TYPE(18)) trunci6(
    .ins (muli2_result),
    .ins_valid (muli2_result_valid),
    .ins_ready (muli2_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci6_outs),
    .outs_valid (trunci6_outs_valid),
    .outs_ready (trunci6_outs_ready)
  );

  oehb #(.DATA_TYPE(14)) buffer56(
    .ins (mux7_outs),
    .ins_valid (mux7_outs_valid),
    .ins_ready (mux7_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer56_outs),
    .outs_valid (buffer56_outs_valid),
    .outs_ready (buffer56_outs_ready)
  );

  tehb #(.DATA_TYPE(14)) buffer57(
    .ins (buffer56_outs),
    .ins_valid (buffer56_outs_valid),
    .ins_ready (buffer56_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer57_outs),
    .outs_valid (buffer57_outs_valid),
    .outs_ready (buffer57_outs_ready)
  );

  extsi #(.INPUT_TYPE(14), .OUTPUT_TYPE(19)) extsi11(
    .ins (buffer57_outs),
    .ins_valid (buffer57_outs_valid),
    .ins_ready (buffer57_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi11_outs),
    .outs_valid (extsi11_outs_valid),
    .outs_ready (extsi11_outs_ready)
  );

  shli #(.DATA_TYPE(19)) shli2(
    .lhs (extsi11_outs),
    .lhs_valid (extsi11_outs_valid),
    .lhs_ready (extsi11_outs_ready),
    .rhs (extsi95_outs),
    .rhs_valid (extsi95_outs_valid),
    .rhs_ready (extsi95_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli2_result),
    .result_valid (shli2_result_valid),
    .result_ready (shli2_result_ready)
  );

  trunci #(.INPUT_TYPE(19), .OUTPUT_TYPE(18)) trunci26(
    .ins (shli2_result),
    .ins_valid (shli2_result_valid),
    .ins_ready (shli2_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci26_outs),
    .outs_valid (trunci26_outs_valid),
    .outs_ready (trunci26_outs_ready)
  );

  addi #(.DATA_TYPE(18)) addi2(
    .lhs (trunci6_outs),
    .lhs_valid (trunci6_outs_valid),
    .lhs_ready (trunci6_outs_ready),
    .rhs (trunci26_outs),
    .rhs_valid (trunci26_outs_valid),
    .rhs_ready (trunci26_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi2_result),
    .result_valid (addi2_result_valid),
    .result_ready (addi2_result_ready)
  );

  extsi #(.INPUT_TYPE(18), .OUTPUT_TYPE(23)) extsi157(
    .ins (addi2_result),
    .ins_valid (addi2_result_valid),
    .ins_ready (addi2_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi157_outs),
    .outs_valid (extsi157_outs_valid),
    .outs_ready (extsi157_outs_ready)
  );

  muli #(.DATA_TYPE(23)) muli3(
    .lhs (extsi157_outs),
    .lhs_valid (extsi157_outs_valid),
    .lhs_ready (extsi157_outs_ready),
    .rhs (extsi148_outs),
    .rhs_valid (extsi148_outs_valid),
    .rhs_ready (extsi148_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli3_result),
    .result_valid (muli3_result_valid),
    .result_ready (muli3_result_ready)
  );

  trunci #(.INPUT_TYPE(23), .OUTPUT_TYPE(21)) trunci8(
    .ins (muli3_result),
    .ins_valid (muli3_result_valid),
    .ins_ready (muli3_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci8_outs),
    .outs_valid (trunci8_outs_valid),
    .outs_ready (trunci8_outs_ready)
  );

  oehb #(.DATA_TYPE(18)) buffer54(
    .ins (mux6_outs),
    .ins_valid (mux6_outs_valid),
    .ins_ready (mux6_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer54_outs),
    .outs_valid (buffer54_outs_valid),
    .outs_ready (buffer54_outs_ready)
  );

  tehb #(.DATA_TYPE(18)) buffer55(
    .ins (buffer54_outs),
    .ins_valid (buffer54_outs_valid),
    .ins_ready (buffer54_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer55_outs),
    .outs_valid (buffer55_outs_valid),
    .outs_ready (buffer55_outs_ready)
  );

  extsi #(.INPUT_TYPE(18), .OUTPUT_TYPE(22)) extsi15(
    .ins (buffer55_outs),
    .ins_valid (buffer55_outs_valid),
    .ins_ready (buffer55_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi15_outs),
    .outs_valid (extsi15_outs_valid),
    .outs_ready (extsi15_outs_ready)
  );

  shli #(.DATA_TYPE(22)) shli3(
    .lhs (extsi15_outs),
    .lhs_valid (extsi15_outs_valid),
    .lhs_ready (extsi15_outs_ready),
    .rhs (extsi94_outs),
    .rhs_valid (extsi94_outs_valid),
    .rhs_ready (extsi94_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli3_result),
    .result_valid (shli3_result_valid),
    .result_ready (shli3_result_ready)
  );

  trunci #(.INPUT_TYPE(22), .OUTPUT_TYPE(21)) trunci27(
    .ins (shli3_result),
    .ins_valid (shli3_result_valid),
    .ins_ready (shli3_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci27_outs),
    .outs_valid (trunci27_outs_valid),
    .outs_ready (trunci27_outs_ready)
  );

  addi #(.DATA_TYPE(21)) addi3(
    .lhs (trunci8_outs),
    .lhs_valid (trunci8_outs_valid),
    .lhs_ready (trunci8_outs_ready),
    .rhs (trunci27_outs),
    .rhs_valid (trunci27_outs_valid),
    .rhs_ready (trunci27_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi3_result),
    .result_valid (addi3_result_valid),
    .result_ready (addi3_result_ready)
  );

  extsi #(.INPUT_TYPE(21), .OUTPUT_TYPE(26)) extsi158(
    .ins (addi3_result),
    .ins_valid (addi3_result_valid),
    .ins_ready (addi3_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi158_outs),
    .outs_valid (extsi158_outs_valid),
    .outs_ready (extsi158_outs_ready)
  );

  muli #(.DATA_TYPE(26)) muli4(
    .lhs (extsi158_outs),
    .lhs_valid (extsi158_outs_valid),
    .lhs_ready (extsi158_outs_ready),
    .rhs (extsi149_outs),
    .rhs_valid (extsi149_outs_valid),
    .rhs_ready (extsi149_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli4_result),
    .result_valid (muli4_result_valid),
    .result_ready (muli4_result_ready)
  );

  trunci #(.INPUT_TYPE(26), .OUTPUT_TYPE(24)) trunci10(
    .ins (muli4_result),
    .ins_valid (muli4_result_valid),
    .ins_ready (muli4_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci10_outs),
    .outs_valid (trunci10_outs_valid),
    .outs_ready (trunci10_outs_ready)
  );

  oehb #(.DATA_TYPE(21)) buffer52(
    .ins (mux5_outs),
    .ins_valid (mux5_outs_valid),
    .ins_ready (mux5_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer52_outs),
    .outs_valid (buffer52_outs_valid),
    .outs_ready (buffer52_outs_ready)
  );

  tehb #(.DATA_TYPE(21)) buffer53(
    .ins (buffer52_outs),
    .ins_valid (buffer52_outs_valid),
    .ins_ready (buffer52_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer53_outs),
    .outs_valid (buffer53_outs_valid),
    .outs_ready (buffer53_outs_ready)
  );

  extsi #(.INPUT_TYPE(21), .OUTPUT_TYPE(25)) extsi19(
    .ins (buffer53_outs),
    .ins_valid (buffer53_outs_valid),
    .ins_ready (buffer53_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi19_outs),
    .outs_valid (extsi19_outs_valid),
    .outs_ready (extsi19_outs_ready)
  );

  shli #(.DATA_TYPE(25)) shli4(
    .lhs (extsi19_outs),
    .lhs_valid (extsi19_outs_valid),
    .lhs_ready (extsi19_outs_ready),
    .rhs (extsi93_outs),
    .rhs_valid (extsi93_outs_valid),
    .rhs_ready (extsi93_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli4_result),
    .result_valid (shli4_result_valid),
    .result_ready (shli4_result_ready)
  );

  trunci #(.INPUT_TYPE(25), .OUTPUT_TYPE(24)) trunci28(
    .ins (shli4_result),
    .ins_valid (shli4_result_valid),
    .ins_ready (shli4_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci28_outs),
    .outs_valid (trunci28_outs_valid),
    .outs_ready (trunci28_outs_ready)
  );

  addi #(.DATA_TYPE(24)) addi4(
    .lhs (trunci10_outs),
    .lhs_valid (trunci10_outs_valid),
    .lhs_ready (trunci10_outs_ready),
    .rhs (trunci28_outs),
    .rhs_valid (trunci28_outs_valid),
    .rhs_ready (trunci28_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi4_result),
    .result_valid (addi4_result_valid),
    .result_ready (addi4_result_ready)
  );

  extsi #(.INPUT_TYPE(24), .OUTPUT_TYPE(29)) extsi159(
    .ins (addi4_result),
    .ins_valid (addi4_result_valid),
    .ins_ready (addi4_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi159_outs),
    .outs_valid (extsi159_outs_valid),
    .outs_ready (extsi159_outs_ready)
  );

  muli #(.DATA_TYPE(29)) muli5(
    .lhs (extsi159_outs),
    .lhs_valid (extsi159_outs_valid),
    .lhs_ready (extsi159_outs_ready),
    .rhs (extsi150_outs),
    .rhs_valid (extsi150_outs_valid),
    .rhs_ready (extsi150_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli5_result),
    .result_valid (muli5_result_valid),
    .result_ready (muli5_result_ready)
  );

  trunci #(.INPUT_TYPE(29), .OUTPUT_TYPE(27)) trunci12(
    .ins (muli5_result),
    .ins_valid (muli5_result_valid),
    .ins_ready (muli5_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci12_outs),
    .outs_valid (trunci12_outs_valid),
    .outs_ready (trunci12_outs_ready)
  );

  oehb #(.DATA_TYPE(24)) buffer50(
    .ins (mux4_outs),
    .ins_valid (mux4_outs_valid),
    .ins_ready (mux4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer50_outs),
    .outs_valid (buffer50_outs_valid),
    .outs_ready (buffer50_outs_ready)
  );

  tehb #(.DATA_TYPE(24)) buffer51(
    .ins (buffer50_outs),
    .ins_valid (buffer50_outs_valid),
    .ins_ready (buffer50_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer51_outs),
    .outs_valid (buffer51_outs_valid),
    .outs_ready (buffer51_outs_ready)
  );

  extsi #(.INPUT_TYPE(24), .OUTPUT_TYPE(28)) extsi23(
    .ins (buffer51_outs),
    .ins_valid (buffer51_outs_valid),
    .ins_ready (buffer51_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi23_outs),
    .outs_valid (extsi23_outs_valid),
    .outs_ready (extsi23_outs_ready)
  );

  shli #(.DATA_TYPE(28)) shli5(
    .lhs (extsi23_outs),
    .lhs_valid (extsi23_outs_valid),
    .lhs_ready (extsi23_outs_ready),
    .rhs (extsi92_outs),
    .rhs_valid (extsi92_outs_valid),
    .rhs_ready (extsi92_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli5_result),
    .result_valid (shli5_result_valid),
    .result_ready (shli5_result_ready)
  );

  trunci #(.INPUT_TYPE(28), .OUTPUT_TYPE(27)) trunci29(
    .ins (shli5_result),
    .ins_valid (shli5_result_valid),
    .ins_ready (shli5_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci29_outs),
    .outs_valid (trunci29_outs_valid),
    .outs_ready (trunci29_outs_ready)
  );

  addi #(.DATA_TYPE(27)) addi5(
    .lhs (trunci12_outs),
    .lhs_valid (trunci12_outs_valid),
    .lhs_ready (trunci12_outs_ready),
    .rhs (trunci29_outs),
    .rhs_valid (trunci29_outs_valid),
    .rhs_ready (trunci29_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi5_result),
    .result_valid (addi5_result_valid),
    .result_ready (addi5_result_ready)
  );

  extsi #(.INPUT_TYPE(27), .OUTPUT_TYPE(32)) extsi160(
    .ins (addi5_result),
    .ins_valid (addi5_result_valid),
    .ins_ready (addi5_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi160_outs),
    .outs_valid (extsi160_outs_valid),
    .outs_ready (extsi160_outs_ready)
  );

  muli #(.DATA_TYPE(32)) muli6(
    .lhs (extsi160_outs),
    .lhs_valid (extsi160_outs_valid),
    .lhs_ready (extsi160_outs_ready),
    .rhs (extsi151_outs),
    .rhs_valid (extsi151_outs_valid),
    .rhs_ready (extsi151_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli6_result),
    .result_valid (muli6_result_valid),
    .result_ready (muli6_result_ready)
  );

  trunci #(.INPUT_TYPE(32), .OUTPUT_TYPE(30)) trunci14(
    .ins (muli6_result),
    .ins_valid (muli6_result_valid),
    .ins_ready (muli6_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci14_outs),
    .outs_valid (trunci14_outs_valid),
    .outs_ready (trunci14_outs_ready)
  );

  oehb #(.DATA_TYPE(27)) buffer48(
    .ins (mux3_outs),
    .ins_valid (mux3_outs_valid),
    .ins_ready (mux3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer48_outs),
    .outs_valid (buffer48_outs_valid),
    .outs_ready (buffer48_outs_ready)
  );

  tehb #(.DATA_TYPE(27)) buffer49(
    .ins (buffer48_outs),
    .ins_valid (buffer48_outs_valid),
    .ins_ready (buffer48_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer49_outs),
    .outs_valid (buffer49_outs_valid),
    .outs_ready (buffer49_outs_ready)
  );

  extsi #(.INPUT_TYPE(27), .OUTPUT_TYPE(31)) extsi27(
    .ins (buffer49_outs),
    .ins_valid (buffer49_outs_valid),
    .ins_ready (buffer49_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi27_outs),
    .outs_valid (extsi27_outs_valid),
    .outs_ready (extsi27_outs_ready)
  );

  shli #(.DATA_TYPE(31)) shli6(
    .lhs (extsi27_outs),
    .lhs_valid (extsi27_outs_valid),
    .lhs_ready (extsi27_outs_ready),
    .rhs (extsi91_outs),
    .rhs_valid (extsi91_outs_valid),
    .rhs_ready (extsi91_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli6_result),
    .result_valid (shli6_result_valid),
    .result_ready (shli6_result_ready)
  );

  trunci #(.INPUT_TYPE(31), .OUTPUT_TYPE(30)) trunci30(
    .ins (shli6_result),
    .ins_valid (shli6_result_valid),
    .ins_ready (shli6_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci30_outs),
    .outs_valid (trunci30_outs_valid),
    .outs_ready (trunci30_outs_ready)
  );

  addi #(.DATA_TYPE(30)) addi6(
    .lhs (trunci14_outs),
    .lhs_valid (trunci14_outs_valid),
    .lhs_ready (trunci14_outs_ready),
    .rhs (trunci30_outs),
    .rhs_valid (trunci30_outs_valid),
    .rhs_ready (trunci30_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi6_result),
    .result_valid (addi6_result_valid),
    .result_ready (addi6_result_ready)
  );

  extsi #(.INPUT_TYPE(30), .OUTPUT_TYPE(35)) extsi161(
    .ins (addi6_result),
    .ins_valid (addi6_result_valid),
    .ins_ready (addi6_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi161_outs),
    .outs_valid (extsi161_outs_valid),
    .outs_ready (extsi161_outs_ready)
  );

  muli #(.DATA_TYPE(35)) muli7(
    .lhs (extsi161_outs),
    .lhs_valid (extsi161_outs_valid),
    .lhs_ready (extsi161_outs_ready),
    .rhs (extsi152_outs),
    .rhs_valid (extsi152_outs_valid),
    .rhs_ready (extsi152_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli7_result),
    .result_valid (muli7_result_valid),
    .result_ready (muli7_result_ready)
  );

  trunci #(.INPUT_TYPE(35), .OUTPUT_TYPE(33)) trunci16(
    .ins (muli7_result),
    .ins_valid (muli7_result_valid),
    .ins_ready (muli7_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci16_outs),
    .outs_valid (trunci16_outs_valid),
    .outs_ready (trunci16_outs_ready)
  );

  oehb #(.DATA_TYPE(30)) buffer46(
    .ins (mux2_outs),
    .ins_valid (mux2_outs_valid),
    .ins_ready (mux2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer46_outs),
    .outs_valid (buffer46_outs_valid),
    .outs_ready (buffer46_outs_ready)
  );

  tehb #(.DATA_TYPE(30)) buffer47(
    .ins (buffer46_outs),
    .ins_valid (buffer46_outs_valid),
    .ins_ready (buffer46_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer47_outs),
    .outs_valid (buffer47_outs_valid),
    .outs_ready (buffer47_outs_ready)
  );

  extsi #(.INPUT_TYPE(30), .OUTPUT_TYPE(34)) extsi31(
    .ins (buffer47_outs),
    .ins_valid (buffer47_outs_valid),
    .ins_ready (buffer47_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi31_outs),
    .outs_valid (extsi31_outs_valid),
    .outs_ready (extsi31_outs_ready)
  );

  shli #(.DATA_TYPE(34)) shli7(
    .lhs (extsi31_outs),
    .lhs_valid (extsi31_outs_valid),
    .lhs_ready (extsi31_outs_ready),
    .rhs (extsi90_outs),
    .rhs_valid (extsi90_outs_valid),
    .rhs_ready (extsi90_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli7_result),
    .result_valid (shli7_result_valid),
    .result_ready (shli7_result_ready)
  );

  trunci #(.INPUT_TYPE(34), .OUTPUT_TYPE(33)) trunci31(
    .ins (shli7_result),
    .ins_valid (shli7_result_valid),
    .ins_ready (shli7_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci31_outs),
    .outs_valid (trunci31_outs_valid),
    .outs_ready (trunci31_outs_ready)
  );

  addi #(.DATA_TYPE(33)) addi7(
    .lhs (trunci16_outs),
    .lhs_valid (trunci16_outs_valid),
    .lhs_ready (trunci16_outs_ready),
    .rhs (trunci31_outs),
    .rhs_valid (trunci31_outs_valid),
    .rhs_ready (trunci31_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi7_result),
    .result_valid (addi7_result_valid),
    .result_ready (addi7_result_ready)
  );

  extsi #(.INPUT_TYPE(33), .OUTPUT_TYPE(38)) extsi162(
    .ins (addi7_result),
    .ins_valid (addi7_result_valid),
    .ins_ready (addi7_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi162_outs),
    .outs_valid (extsi162_outs_valid),
    .outs_ready (extsi162_outs_ready)
  );

  muli #(.DATA_TYPE(38)) muli8(
    .lhs (extsi162_outs),
    .lhs_valid (extsi162_outs_valid),
    .lhs_ready (extsi162_outs_ready),
    .rhs (extsi153_outs),
    .rhs_valid (extsi153_outs_valid),
    .rhs_ready (extsi153_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli8_result),
    .result_valid (muli8_result_valid),
    .result_ready (muli8_result_ready)
  );

  trunci #(.INPUT_TYPE(38), .OUTPUT_TYPE(37)) trunci18(
    .ins (muli8_result),
    .ins_valid (muli8_result_valid),
    .ins_ready (muli8_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci18_outs),
    .outs_valid (trunci18_outs_valid),
    .outs_ready (trunci18_outs_ready)
  );

  oehb #(.DATA_TYPE(34)) buffer44(
    .ins (mux1_outs),
    .ins_valid (mux1_outs_valid),
    .ins_ready (mux1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer44_outs),
    .outs_valid (buffer44_outs_valid),
    .outs_ready (buffer44_outs_ready)
  );

  tehb #(.DATA_TYPE(34)) buffer45(
    .ins (buffer44_outs),
    .ins_valid (buffer44_outs_valid),
    .ins_ready (buffer44_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer45_outs),
    .outs_valid (buffer45_outs_valid),
    .outs_ready (buffer45_outs_ready)
  );

  extsi #(.INPUT_TYPE(34), .OUTPUT_TYPE(38)) extsi35(
    .ins (buffer45_outs),
    .ins_valid (buffer45_outs_valid),
    .ins_ready (buffer45_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi35_outs),
    .outs_valid (extsi35_outs_valid),
    .outs_ready (extsi35_outs_ready)
  );

  shli #(.DATA_TYPE(38)) shli8(
    .lhs (extsi35_outs),
    .lhs_valid (extsi35_outs_valid),
    .lhs_ready (extsi35_outs_ready),
    .rhs (extsi89_outs),
    .rhs_valid (extsi89_outs_valid),
    .rhs_ready (extsi89_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli8_result),
    .result_valid (shli8_result_valid),
    .result_ready (shli8_result_ready)
  );

  trunci #(.INPUT_TYPE(38), .OUTPUT_TYPE(37)) trunci32(
    .ins (shli8_result),
    .ins_valid (shli8_result_valid),
    .ins_ready (shli8_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci32_outs),
    .outs_valid (trunci32_outs_valid),
    .outs_ready (trunci32_outs_ready)
  );

  addi #(.DATA_TYPE(37)) addi8(
    .lhs (trunci18_outs),
    .lhs_valid (trunci18_outs_valid),
    .lhs_ready (trunci18_outs_ready),
    .rhs (trunci32_outs),
    .rhs_valid (trunci32_outs_valid),
    .rhs_ready (trunci32_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi8_result),
    .result_valid (addi8_result_valid),
    .result_ready (addi8_result_ready)
  );

  extsi #(.INPUT_TYPE(37), .OUTPUT_TYPE(42)) extsi163(
    .ins (addi8_result),
    .ins_valid (addi8_result_valid),
    .ins_ready (addi8_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi163_outs),
    .outs_valid (extsi163_outs_valid),
    .outs_ready (extsi163_outs_ready)
  );

  muli #(.DATA_TYPE(42)) muli9(
    .lhs (extsi163_outs),
    .lhs_valid (extsi163_outs_valid),
    .lhs_ready (extsi163_outs_ready),
    .rhs (extsi154_outs),
    .rhs_valid (extsi154_outs_valid),
    .rhs_ready (extsi154_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli9_result),
    .result_valid (muli9_result_valid),
    .result_ready (muli9_result_ready)
  );

  trunci #(.INPUT_TYPE(42), .OUTPUT_TYPE(13)) trunci33(
    .ins (muli9_result),
    .ins_valid (muli9_result_valid),
    .ins_ready (muli9_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci33_outs),
    .outs_valid (trunci33_outs_valid),
    .outs_ready (trunci33_outs_ready)
  );

  oehb #(.DATA_TYPE(36)) buffer42(
    .ins (mux0_outs),
    .ins_valid (mux0_outs_valid),
    .ins_ready (mux0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer42_outs),
    .outs_valid (buffer42_outs_valid),
    .outs_ready (buffer42_outs_ready)
  );

  tehb #(.DATA_TYPE(36)) buffer43(
    .ins (buffer42_outs),
    .ins_valid (buffer42_outs_valid),
    .ins_ready (buffer42_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer43_outs),
    .outs_valid (buffer43_outs_valid),
    .outs_ready (buffer43_outs_ready)
  );

  extsi #(.INPUT_TYPE(36), .OUTPUT_TYPE(40)) extsi39(
    .ins (buffer43_outs),
    .ins_valid (buffer43_outs_valid),
    .ins_ready (buffer43_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi39_outs),
    .outs_valid (extsi39_outs_valid),
    .outs_ready (extsi39_outs_ready)
  );

  shli #(.DATA_TYPE(40)) shli9(
    .lhs (extsi39_outs),
    .lhs_valid (extsi39_outs_valid),
    .lhs_ready (extsi39_outs_ready),
    .rhs (extsi88_outs),
    .rhs_valid (extsi88_outs_valid),
    .rhs_ready (extsi88_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli9_result),
    .result_valid (shli9_result_valid),
    .result_ready (shli9_result_ready)
  );

  trunci #(.INPUT_TYPE(40), .OUTPUT_TYPE(13)) trunci34(
    .ins (shli9_result),
    .ins_valid (shli9_result_valid),
    .ins_ready (shli9_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci34_outs),
    .outs_valid (trunci34_outs_valid),
    .outs_ready (trunci34_outs_ready)
  );

  addi #(.DATA_TYPE(13)) addi9(
    .lhs (trunci33_outs),
    .lhs_valid (trunci33_outs_valid),
    .lhs_ready (trunci33_outs_ready),
    .rhs (trunci34_outs),
    .rhs_valid (trunci34_outs_valid),
    .rhs_ready (trunci34_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi9_result),
    .result_valid (addi9_result_valid),
    .result_ready (addi9_result_ready)
  );

  shrsi #(.DATA_TYPE(13)) shrsi0(
    .lhs (addi9_result),
    .lhs_valid (addi9_result_valid),
    .lhs_ready (addi9_result_ready),
    .rhs (extui0_outs),
    .rhs_valid (extui0_outs_valid),
    .rhs_ready (extui0_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shrsi0_result),
    .result_valid (shrsi0_result_valid),
    .result_ready (shrsi0_result_ready)
  );

  trunci #(.INPUT_TYPE(13), .OUTPUT_TYPE(8)) trunci22(
    .ins (shrsi0_result),
    .ins_valid (shrsi0_result_valid),
    .ins_ready (shrsi0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci22_outs),
    .outs_valid (trunci22_outs_valid),
    .outs_ready (trunci22_outs_ready)
  );

endmodule
