/*
 * Copyright (c) 2024 Louis Ledoux, Pierre Cochard, Emeraude Team @INRIA
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module ttgf0p2_faust_top (
    input  wire [7:0] ui_in,    // Dedicated inputs (unused here)
    output wire [7:0] uo_out,   // Dedicated outputs -> R-2R ladder
    input  wire [7:0] uio_in,   // Bidirectional IOs: input path
    output wire [7:0] uio_out,  // Bidirectional IOs: output path
    output wire [7:0] uio_oe,   // Bidirectional IOs: output enable (1=output)
    input  wire       ena,      // Always 1 when powered
    input  wire       clk,      // Global clock
    input  wire       rst_n     // Active-low reset
);

  // ---------------------------------------------------------------------------
  // Internal wires
  // ---------------------------------------------------------------------------
  wire [15:0] faust_sample;   // Full-precision sample from Faust
  wire [7:0]  audio_out;      // Truncated 8-bit sample for DAC

  // ---------------------------------------------------------------------------
  // Faust DSP core instance
  // ---------------------------------------------------------------------------
  // The core should output one sample per clock
  faust_core core (
      .clk  (clk),
      .rst  (!rst_n),          // Convert active-low reset to active-high
      .out  (faust_sample)     // 16-bit signed or unsigned output
  );

  // ---------------------------------------------------------------------------
  // Output truncation / quantization
  // TODO: check what outputs faust
  // ---------------------------------------------------------------------------
  assign audio_out = faust_sample[15:8];  // Simple 8-bit truncation
  assign uo_out    = audio_out;           // Drive R-2R DAC outputs

  // ---------------------------------------------------------------------------
  // Unused IO configuration
  // ---------------------------------------------------------------------------
  assign uio_out = 8'b0;   // Not used
  assign uio_oe  = 8'b0;   // Configure all UIO pins as inputs

  // Tie off unused inputs to prevent synthesis warnings
  wire _unused = &{ena, ui_in, uio_in, 1'b0};

endmodule