module process(
  input [16:0] in0,
  input  in0_valid,
  input  start_valid,
  input  clk,
  input  rst,
  input  out0_ready,
  input  end_ready,
  output  in0_ready,
  output  start_ready,
  output [7:0] out0,
  output  out0_valid,
  output  end_valid
);
  wire  fork0_outs_0_valid;
  wire  fork0_outs_0_ready;
  wire  fork0_outs_1_valid;
  wire  fork0_outs_1_ready;
  wire  fork0_outs_2_valid;
  wire  fork0_outs_2_ready;
  wire  fork0_outs_3_valid;
  wire  fork0_outs_3_ready;
  wire  fork0_outs_4_valid;
  wire  fork0_outs_4_ready;
  wire  fork0_outs_5_valid;
  wire  fork0_outs_5_ready;
  wire  fork0_outs_6_valid;
  wire  fork0_outs_6_ready;
  wire  fork0_outs_7_valid;
  wire  fork0_outs_7_ready;
  wire [16:0] fork1_outs_0;
  wire  fork1_outs_0_valid;
  wire  fork1_outs_0_ready;
  wire [16:0] fork1_outs_1;
  wire  fork1_outs_1_valid;
  wire  fork1_outs_1_ready;
  wire [6:0] trunci13_outs;
  wire  trunci13_outs_valid;
  wire  trunci13_outs_ready;
  wire  source0_outs_valid;
  wire  source0_outs_ready;
  wire [0:0] constant459_outs;
  wire  constant459_outs_valid;
  wire  constant459_outs_ready;
  wire [4:0] extsi141_outs;
  wire  extsi141_outs_valid;
  wire  extsi141_outs_ready;
  wire [11:0] constant223_outs;
  wire  constant223_outs_valid;
  wire  constant223_outs_ready;
  wire [14:0] constant460_outs;
  wire  constant460_outs_valid;
  wire  constant460_outs_ready;
  wire [21:0] constant225_outs;
  wire  constant225_outs_valid;
  wire  constant225_outs_ready;
  wire [26:0] constant226_outs;
  wire  constant226_outs_valid;
  wire  constant226_outs_ready;
  wire [32:0] constant227_outs;
  wire  constant227_outs_valid;
  wire  constant227_outs_ready;
  wire [32:0] constant461_outs;
  wire  constant461_outs_valid;
  wire  constant461_outs_ready;
  wire  source1_outs_valid;
  wire  source1_outs_ready;
  wire [4:0] constant462_outs;
  wire  constant462_outs_valid;
  wire  constant462_outs_ready;
  wire [16:0] extsi23_outs;
  wire  extsi23_outs_valid;
  wire  extsi23_outs_ready;
  wire [16:0] shrui0_result;
  wire  shrui0_result_valid;
  wire  shrui0_result_ready;
  wire [4:0] trunci0_outs;
  wire  trunci0_outs_valid;
  wire  trunci0_outs_ready;
  wire [4:0] fork2_outs_0;
  wire  fork2_outs_0_valid;
  wire  fork2_outs_0_ready;
  wire [4:0] fork2_outs_1;
  wire  fork2_outs_1_valid;
  wire  fork2_outs_1_ready;
  wire [0:0] cmpi0_result;
  wire  cmpi0_result_valid;
  wire  cmpi0_result_ready;
  wire [0:0] fork3_outs_0;
  wire  fork3_outs_0_valid;
  wire  fork3_outs_0_ready;
  wire [0:0] fork3_outs_1;
  wire  fork3_outs_1_valid;
  wire  fork3_outs_1_ready;
  wire [0:0] fork3_outs_2;
  wire  fork3_outs_2_valid;
  wire  fork3_outs_2_ready;
  wire [0:0] fork3_outs_3;
  wire  fork3_outs_3_valid;
  wire  fork3_outs_3_ready;
  wire [0:0] fork3_outs_4;
  wire  fork3_outs_4_valid;
  wire  fork3_outs_4_ready;
  wire [0:0] fork3_outs_5;
  wire  fork3_outs_5_valid;
  wire  fork3_outs_5_ready;
  wire [0:0] fork3_outs_6;
  wire  fork3_outs_6_valid;
  wire  fork3_outs_6_ready;
  wire [0:0] fork3_outs_7;
  wire  fork3_outs_7_valid;
  wire  fork3_outs_7_ready;
  wire [0:0] fork3_outs_8;
  wire  fork3_outs_8_valid;
  wire  fork3_outs_8_ready;
  wire [32:0] cond_br32_trueOut;
  wire  cond_br32_trueOut_valid;
  wire  cond_br32_trueOut_ready;
  wire [32:0] cond_br32_falseOut;
  wire  cond_br32_falseOut_valid;
  wire  cond_br32_falseOut_ready;
  wire [36:0] extsi142_outs;
  wire  extsi142_outs_valid;
  wire  extsi142_outs_ready;
  wire [32:0] cond_br33_trueOut;
  wire  cond_br33_trueOut_valid;
  wire  cond_br33_trueOut_ready;
  wire [32:0] cond_br33_falseOut;
  wire  cond_br33_falseOut_valid;
  wire  cond_br33_falseOut_ready;
  wire [26:0] cond_br34_trueOut;
  wire  cond_br34_trueOut_valid;
  wire  cond_br34_trueOut_ready;
  wire [26:0] cond_br34_falseOut;
  wire  cond_br34_falseOut_valid;
  wire  cond_br34_falseOut_ready;
  wire [21:0] cond_br35_trueOut;
  wire  cond_br35_trueOut_valid;
  wire  cond_br35_trueOut_ready;
  wire [21:0] cond_br35_falseOut;
  wire  cond_br35_falseOut_valid;
  wire  cond_br35_falseOut_ready;
  wire [14:0] cond_br36_trueOut;
  wire  cond_br36_trueOut_valid;
  wire  cond_br36_trueOut_ready;
  wire [14:0] cond_br36_falseOut;
  wire  cond_br36_falseOut_valid;
  wire  cond_br36_falseOut_ready;
  wire [16:0] extsi143_outs;
  wire  extsi143_outs_valid;
  wire  extsi143_outs_ready;
  wire [11:0] cond_br37_trueOut;
  wire  cond_br37_trueOut_valid;
  wire  cond_br37_trueOut_ready;
  wire [11:0] cond_br37_falseOut;
  wire  cond_br37_falseOut_valid;
  wire  cond_br37_falseOut_ready;
  wire [6:0] cond_br38_trueOut;
  wire  cond_br38_trueOut_valid;
  wire  cond_br38_trueOut_ready;
  wire [6:0] cond_br38_falseOut;
  wire  cond_br38_falseOut_valid;
  wire  cond_br38_falseOut_ready;
  wire  cond_br39_trueOut_valid;
  wire  cond_br39_trueOut_ready;
  wire  cond_br39_falseOut_valid;
  wire  cond_br39_falseOut_ready;
  wire [4:0] cond_br40_trueOut;
  wire  cond_br40_trueOut_valid;
  wire  cond_br40_trueOut_ready;
  wire [4:0] cond_br40_falseOut;
  wire  cond_br40_falseOut_valid;
  wire  cond_br40_falseOut_ready;
  wire [4:0] buffer2_outs;
  wire  buffer2_outs_valid;
  wire  buffer2_outs_ready;
  wire [4:0] buffer3_outs;
  wire  buffer3_outs_valid;
  wire  buffer3_outs_ready;
  wire [4:0] fork4_outs_0;
  wire  fork4_outs_0_valid;
  wire  fork4_outs_0_ready;
  wire [4:0] fork4_outs_1;
  wire  fork4_outs_1_valid;
  wire  fork4_outs_1_ready;
  wire  buffer4_outs_valid;
  wire  buffer4_outs_ready;
  wire  buffer5_outs_valid;
  wire  buffer5_outs_ready;
  wire  fork5_outs_0_valid;
  wire  fork5_outs_0_ready;
  wire  fork5_outs_1_valid;
  wire  fork5_outs_1_ready;
  wire  fork5_outs_2_valid;
  wire  fork5_outs_2_ready;
  wire  fork5_outs_3_valid;
  wire  fork5_outs_3_ready;
  wire  fork5_outs_4_valid;
  wire  fork5_outs_4_ready;
  wire  fork5_outs_5_valid;
  wire  fork5_outs_5_ready;
  wire  fork5_outs_6_valid;
  wire  fork5_outs_6_ready;
  wire [33:0] constant463_outs;
  wire  constant463_outs_valid;
  wire  constant463_outs_ready;
  wire [32:0] constant231_outs;
  wire  constant231_outs_valid;
  wire  constant231_outs_ready;
  wire [26:0] constant232_outs;
  wire  constant232_outs_valid;
  wire  constant232_outs_ready;
  wire [21:0] constant233_outs;
  wire  constant233_outs_valid;
  wire  constant233_outs_ready;
  wire [15:0] constant464_outs;
  wire  constant464_outs_valid;
  wire  constant464_outs_ready;
  wire [11:0] constant235_outs;
  wire  constant235_outs_valid;
  wire  constant235_outs_ready;
  wire  source2_outs_valid;
  wire  source2_outs_ready;
  wire [1:0] constant465_outs;
  wire  constant465_outs_valid;
  wire  constant465_outs_ready;
  wire [4:0] extsi144_outs;
  wire  extsi144_outs_valid;
  wire  extsi144_outs_ready;
  wire [0:0] cmpi1_result;
  wire  cmpi1_result_valid;
  wire  cmpi1_result_ready;
  wire [0:0] fork6_outs_0;
  wire  fork6_outs_0_valid;
  wire  fork6_outs_0_ready;
  wire [0:0] fork6_outs_1;
  wire  fork6_outs_1_valid;
  wire  fork6_outs_1_ready;
  wire [0:0] fork6_outs_2;
  wire  fork6_outs_2_valid;
  wire  fork6_outs_2_ready;
  wire [0:0] fork6_outs_3;
  wire  fork6_outs_3_valid;
  wire  fork6_outs_3_ready;
  wire [0:0] fork6_outs_4;
  wire  fork6_outs_4_valid;
  wire  fork6_outs_4_ready;
  wire [0:0] fork6_outs_5;
  wire  fork6_outs_5_valid;
  wire  fork6_outs_5_ready;
  wire [0:0] fork6_outs_6;
  wire  fork6_outs_6_valid;
  wire  fork6_outs_6_ready;
  wire [0:0] fork6_outs_7;
  wire  fork6_outs_7_valid;
  wire  fork6_outs_7_ready;
  wire [0:0] fork6_outs_8;
  wire  fork6_outs_8_valid;
  wire  fork6_outs_8_ready;
  wire [33:0] cond_br41_trueOut;
  wire  cond_br41_trueOut_valid;
  wire  cond_br41_trueOut_ready;
  wire [33:0] cond_br41_falseOut;
  wire  cond_br41_falseOut_valid;
  wire  cond_br41_falseOut_ready;
  wire [36:0] extsi145_outs;
  wire  extsi145_outs_valid;
  wire  extsi145_outs_ready;
  wire [32:0] cond_br42_trueOut;
  wire  cond_br42_trueOut_valid;
  wire  cond_br42_trueOut_ready;
  wire [32:0] cond_br42_falseOut;
  wire  cond_br42_falseOut_valid;
  wire  cond_br42_falseOut_ready;
  wire [26:0] cond_br43_trueOut;
  wire  cond_br43_trueOut_valid;
  wire  cond_br43_trueOut_ready;
  wire [26:0] cond_br43_falseOut;
  wire  cond_br43_falseOut_valid;
  wire  cond_br43_falseOut_ready;
  wire [21:0] cond_br44_trueOut;
  wire  cond_br44_trueOut_valid;
  wire  cond_br44_trueOut_ready;
  wire [21:0] cond_br44_falseOut;
  wire  cond_br44_falseOut_valid;
  wire  cond_br44_falseOut_ready;
  wire [15:0] cond_br45_trueOut;
  wire  cond_br45_trueOut_valid;
  wire  cond_br45_trueOut_ready;
  wire [15:0] cond_br45_falseOut;
  wire  cond_br45_falseOut_valid;
  wire  cond_br45_falseOut_ready;
  wire [16:0] extsi146_outs;
  wire  extsi146_outs_valid;
  wire  extsi146_outs_ready;
  wire [11:0] cond_br46_trueOut;
  wire  cond_br46_trueOut_valid;
  wire  cond_br46_trueOut_ready;
  wire [11:0] cond_br46_falseOut;
  wire  cond_br46_falseOut_valid;
  wire  cond_br46_falseOut_ready;
  wire [6:0] buffer0_outs;
  wire  buffer0_outs_valid;
  wire  buffer0_outs_ready;
  wire [6:0] buffer1_outs;
  wire  buffer1_outs_valid;
  wire  buffer1_outs_ready;
  wire [6:0] cond_br47_trueOut;
  wire  cond_br47_trueOut_valid;
  wire  cond_br47_trueOut_ready;
  wire [6:0] cond_br47_falseOut;
  wire  cond_br47_falseOut_valid;
  wire  cond_br47_falseOut_ready;
  wire  cond_br48_trueOut_valid;
  wire  cond_br48_trueOut_ready;
  wire  cond_br48_falseOut_valid;
  wire  cond_br48_falseOut_ready;
  wire [4:0] cond_br49_trueOut;
  wire  cond_br49_trueOut_valid;
  wire  cond_br49_trueOut_ready;
  wire [4:0] cond_br49_falseOut;
  wire  cond_br49_falseOut_valid;
  wire  cond_br49_falseOut_ready;
  wire [4:0] buffer8_outs;
  wire  buffer8_outs_valid;
  wire  buffer8_outs_ready;
  wire [4:0] buffer9_outs;
  wire  buffer9_outs_valid;
  wire  buffer9_outs_ready;
  wire [4:0] fork7_outs_0;
  wire  fork7_outs_0_valid;
  wire  fork7_outs_0_ready;
  wire [4:0] fork7_outs_1;
  wire  fork7_outs_1_valid;
  wire  fork7_outs_1_ready;
  wire  buffer10_outs_valid;
  wire  buffer10_outs_ready;
  wire  buffer11_outs_valid;
  wire  buffer11_outs_ready;
  wire  fork8_outs_0_valid;
  wire  fork8_outs_0_ready;
  wire  fork8_outs_1_valid;
  wire  fork8_outs_1_ready;
  wire  fork8_outs_2_valid;
  wire  fork8_outs_2_ready;
  wire  fork8_outs_3_valid;
  wire  fork8_outs_3_ready;
  wire  fork8_outs_4_valid;
  wire  fork8_outs_4_ready;
  wire  fork8_outs_5_valid;
  wire  fork8_outs_5_ready;
  wire  fork8_outs_6_valid;
  wire  fork8_outs_6_ready;
  wire [34:0] constant466_outs;
  wire  constant466_outs_valid;
  wire  constant466_outs_ready;
  wire [32:0] constant238_outs;
  wire  constant238_outs_valid;
  wire  constant238_outs_ready;
  wire [26:0] constant239_outs;
  wire  constant239_outs_valid;
  wire  constant239_outs_ready;
  wire [21:0] constant240_outs;
  wire  constant240_outs_valid;
  wire  constant240_outs_ready;
  wire [16:0] constant241_outs;
  wire  constant241_outs_valid;
  wire  constant241_outs_ready;
  wire [11:0] constant242_outs;
  wire  constant242_outs_valid;
  wire  constant242_outs_ready;
  wire  source3_outs_valid;
  wire  source3_outs_ready;
  wire [2:0] constant467_outs;
  wire  constant467_outs_valid;
  wire  constant467_outs_ready;
  wire [4:0] extsi147_outs;
  wire  extsi147_outs_valid;
  wire  extsi147_outs_ready;
  wire [0:0] cmpi2_result;
  wire  cmpi2_result_valid;
  wire  cmpi2_result_ready;
  wire [0:0] fork9_outs_0;
  wire  fork9_outs_0_valid;
  wire  fork9_outs_0_ready;
  wire [0:0] fork9_outs_1;
  wire  fork9_outs_1_valid;
  wire  fork9_outs_1_ready;
  wire [0:0] fork9_outs_2;
  wire  fork9_outs_2_valid;
  wire  fork9_outs_2_ready;
  wire [0:0] fork9_outs_3;
  wire  fork9_outs_3_valid;
  wire  fork9_outs_3_ready;
  wire [0:0] fork9_outs_4;
  wire  fork9_outs_4_valid;
  wire  fork9_outs_4_ready;
  wire [0:0] fork9_outs_5;
  wire  fork9_outs_5_valid;
  wire  fork9_outs_5_ready;
  wire [0:0] fork9_outs_6;
  wire  fork9_outs_6_valid;
  wire  fork9_outs_6_ready;
  wire [0:0] fork9_outs_7;
  wire  fork9_outs_7_valid;
  wire  fork9_outs_7_ready;
  wire [0:0] fork9_outs_8;
  wire  fork9_outs_8_valid;
  wire  fork9_outs_8_ready;
  wire [34:0] cond_br50_trueOut;
  wire  cond_br50_trueOut_valid;
  wire  cond_br50_trueOut_ready;
  wire [34:0] cond_br50_falseOut;
  wire  cond_br50_falseOut_valid;
  wire  cond_br50_falseOut_ready;
  wire [36:0] extsi148_outs;
  wire  extsi148_outs_valid;
  wire  extsi148_outs_ready;
  wire [32:0] cond_br51_trueOut;
  wire  cond_br51_trueOut_valid;
  wire  cond_br51_trueOut_ready;
  wire [32:0] cond_br51_falseOut;
  wire  cond_br51_falseOut_valid;
  wire  cond_br51_falseOut_ready;
  wire [26:0] cond_br52_trueOut;
  wire  cond_br52_trueOut_valid;
  wire  cond_br52_trueOut_ready;
  wire [26:0] cond_br52_falseOut;
  wire  cond_br52_falseOut_valid;
  wire  cond_br52_falseOut_ready;
  wire [21:0] cond_br53_trueOut;
  wire  cond_br53_trueOut_valid;
  wire  cond_br53_trueOut_ready;
  wire [21:0] cond_br53_falseOut;
  wire  cond_br53_falseOut_valid;
  wire  cond_br53_falseOut_ready;
  wire [16:0] cond_br54_trueOut;
  wire  cond_br54_trueOut_valid;
  wire  cond_br54_trueOut_ready;
  wire [16:0] cond_br54_falseOut;
  wire  cond_br54_falseOut_valid;
  wire  cond_br54_falseOut_ready;
  wire [11:0] cond_br55_trueOut;
  wire  cond_br55_trueOut_valid;
  wire  cond_br55_trueOut_ready;
  wire [11:0] cond_br55_falseOut;
  wire  cond_br55_falseOut_valid;
  wire  cond_br55_falseOut_ready;
  wire [6:0] buffer6_outs;
  wire  buffer6_outs_valid;
  wire  buffer6_outs_ready;
  wire [6:0] buffer7_outs;
  wire  buffer7_outs_valid;
  wire  buffer7_outs_ready;
  wire [6:0] cond_br56_trueOut;
  wire  cond_br56_trueOut_valid;
  wire  cond_br56_trueOut_ready;
  wire [6:0] cond_br56_falseOut;
  wire  cond_br56_falseOut_valid;
  wire  cond_br56_falseOut_ready;
  wire  cond_br57_trueOut_valid;
  wire  cond_br57_trueOut_ready;
  wire  cond_br57_falseOut_valid;
  wire  cond_br57_falseOut_ready;
  wire [4:0] cond_br58_trueOut;
  wire  cond_br58_trueOut_valid;
  wire  cond_br58_trueOut_ready;
  wire [4:0] cond_br58_falseOut;
  wire  cond_br58_falseOut_valid;
  wire  cond_br58_falseOut_ready;
  wire [4:0] buffer14_outs;
  wire  buffer14_outs_valid;
  wire  buffer14_outs_ready;
  wire [4:0] buffer15_outs;
  wire  buffer15_outs_valid;
  wire  buffer15_outs_ready;
  wire [4:0] fork10_outs_0;
  wire  fork10_outs_0_valid;
  wire  fork10_outs_0_ready;
  wire [4:0] fork10_outs_1;
  wire  fork10_outs_1_valid;
  wire  fork10_outs_1_ready;
  wire  buffer16_outs_valid;
  wire  buffer16_outs_ready;
  wire  buffer17_outs_valid;
  wire  buffer17_outs_ready;
  wire  fork11_outs_0_valid;
  wire  fork11_outs_0_ready;
  wire  fork11_outs_1_valid;
  wire  fork11_outs_1_ready;
  wire  fork11_outs_2_valid;
  wire  fork11_outs_2_ready;
  wire  fork11_outs_3_valid;
  wire  fork11_outs_3_ready;
  wire  fork11_outs_4_valid;
  wire  fork11_outs_4_ready;
  wire  fork11_outs_5_valid;
  wire  fork11_outs_5_ready;
  wire  fork11_outs_6_valid;
  wire  fork11_outs_6_ready;
  wire [35:0] constant468_outs;
  wire  constant468_outs_valid;
  wire  constant468_outs_ready;
  wire [32:0] constant245_outs;
  wire  constant245_outs_valid;
  wire  constant245_outs_ready;
  wire [26:0] constant246_outs;
  wire  constant246_outs_valid;
  wire  constant246_outs_ready;
  wire [21:0] constant247_outs;
  wire  constant247_outs_valid;
  wire  constant247_outs_ready;
  wire [16:0] constant248_outs;
  wire  constant248_outs_valid;
  wire  constant248_outs_ready;
  wire [10:0] constant469_outs;
  wire  constant469_outs_valid;
  wire  constant469_outs_ready;
  wire  source4_outs_valid;
  wire  source4_outs_ready;
  wire [2:0] constant470_outs;
  wire  constant470_outs_valid;
  wire  constant470_outs_ready;
  wire [4:0] extsi149_outs;
  wire  extsi149_outs_valid;
  wire  extsi149_outs_ready;
  wire [0:0] cmpi3_result;
  wire  cmpi3_result_valid;
  wire  cmpi3_result_ready;
  wire [0:0] fork12_outs_0;
  wire  fork12_outs_0_valid;
  wire  fork12_outs_0_ready;
  wire [0:0] fork12_outs_1;
  wire  fork12_outs_1_valid;
  wire  fork12_outs_1_ready;
  wire [0:0] fork12_outs_2;
  wire  fork12_outs_2_valid;
  wire  fork12_outs_2_ready;
  wire [0:0] fork12_outs_3;
  wire  fork12_outs_3_valid;
  wire  fork12_outs_3_ready;
  wire [0:0] fork12_outs_4;
  wire  fork12_outs_4_valid;
  wire  fork12_outs_4_ready;
  wire [0:0] fork12_outs_5;
  wire  fork12_outs_5_valid;
  wire  fork12_outs_5_ready;
  wire [0:0] fork12_outs_6;
  wire  fork12_outs_6_valid;
  wire  fork12_outs_6_ready;
  wire [0:0] fork12_outs_7;
  wire  fork12_outs_7_valid;
  wire  fork12_outs_7_ready;
  wire [0:0] fork12_outs_8;
  wire  fork12_outs_8_valid;
  wire  fork12_outs_8_ready;
  wire [35:0] cond_br59_trueOut;
  wire  cond_br59_trueOut_valid;
  wire  cond_br59_trueOut_ready;
  wire [35:0] cond_br59_falseOut;
  wire  cond_br59_falseOut_valid;
  wire  cond_br59_falseOut_ready;
  wire [36:0] extsi150_outs;
  wire  extsi150_outs_valid;
  wire  extsi150_outs_ready;
  wire [32:0] cond_br60_trueOut;
  wire  cond_br60_trueOut_valid;
  wire  cond_br60_trueOut_ready;
  wire [32:0] cond_br60_falseOut;
  wire  cond_br60_falseOut_valid;
  wire  cond_br60_falseOut_ready;
  wire [26:0] cond_br61_trueOut;
  wire  cond_br61_trueOut_valid;
  wire  cond_br61_trueOut_ready;
  wire [26:0] cond_br61_falseOut;
  wire  cond_br61_falseOut_valid;
  wire  cond_br61_falseOut_ready;
  wire [21:0] cond_br62_trueOut;
  wire  cond_br62_trueOut_valid;
  wire  cond_br62_trueOut_ready;
  wire [21:0] cond_br62_falseOut;
  wire  cond_br62_falseOut_valid;
  wire  cond_br62_falseOut_ready;
  wire [16:0] cond_br63_trueOut;
  wire  cond_br63_trueOut_valid;
  wire  cond_br63_trueOut_ready;
  wire [16:0] cond_br63_falseOut;
  wire  cond_br63_falseOut_valid;
  wire  cond_br63_falseOut_ready;
  wire [10:0] cond_br64_trueOut;
  wire  cond_br64_trueOut_valid;
  wire  cond_br64_trueOut_ready;
  wire [10:0] cond_br64_falseOut;
  wire  cond_br64_falseOut_valid;
  wire  cond_br64_falseOut_ready;
  wire [11:0] extsi151_outs;
  wire  extsi151_outs_valid;
  wire  extsi151_outs_ready;
  wire [6:0] buffer12_outs;
  wire  buffer12_outs_valid;
  wire  buffer12_outs_ready;
  wire [6:0] buffer13_outs;
  wire  buffer13_outs_valid;
  wire  buffer13_outs_ready;
  wire [6:0] cond_br65_trueOut;
  wire  cond_br65_trueOut_valid;
  wire  cond_br65_trueOut_ready;
  wire [6:0] cond_br65_falseOut;
  wire  cond_br65_falseOut_valid;
  wire  cond_br65_falseOut_ready;
  wire  cond_br66_trueOut_valid;
  wire  cond_br66_trueOut_ready;
  wire  cond_br66_falseOut_valid;
  wire  cond_br66_falseOut_ready;
  wire [4:0] cond_br67_trueOut;
  wire  cond_br67_trueOut_valid;
  wire  cond_br67_trueOut_ready;
  wire [4:0] cond_br67_falseOut;
  wire  cond_br67_falseOut_valid;
  wire  cond_br67_falseOut_ready;
  wire [4:0] buffer20_outs;
  wire  buffer20_outs_valid;
  wire  buffer20_outs_ready;
  wire [4:0] buffer21_outs;
  wire  buffer21_outs_valid;
  wire  buffer21_outs_ready;
  wire [4:0] fork13_outs_0;
  wire  fork13_outs_0_valid;
  wire  fork13_outs_0_ready;
  wire [4:0] fork13_outs_1;
  wire  fork13_outs_1_valid;
  wire  fork13_outs_1_ready;
  wire  buffer22_outs_valid;
  wire  buffer22_outs_ready;
  wire  buffer23_outs_valid;
  wire  buffer23_outs_ready;
  wire  fork14_outs_0_valid;
  wire  fork14_outs_0_ready;
  wire  fork14_outs_1_valid;
  wire  fork14_outs_1_ready;
  wire  fork14_outs_2_valid;
  wire  fork14_outs_2_ready;
  wire  fork14_outs_3_valid;
  wire  fork14_outs_3_ready;
  wire  fork14_outs_4_valid;
  wire  fork14_outs_4_ready;
  wire  fork14_outs_5_valid;
  wire  fork14_outs_5_ready;
  wire  fork14_outs_6_valid;
  wire  fork14_outs_6_ready;
  wire [35:0] constant471_outs;
  wire  constant471_outs_valid;
  wire  constant471_outs_ready;
  wire [32:0] constant252_outs;
  wire  constant252_outs_valid;
  wire  constant252_outs_ready;
  wire [26:0] constant253_outs;
  wire  constant253_outs_valid;
  wire  constant253_outs_ready;
  wire [21:0] constant254_outs;
  wire  constant254_outs_valid;
  wire  constant254_outs_ready;
  wire [16:0] constant255_outs;
  wire  constant255_outs_valid;
  wire  constant255_outs_ready;
  wire [11:0] constant256_outs;
  wire  constant256_outs_valid;
  wire  constant256_outs_ready;
  wire  source5_outs_valid;
  wire  source5_outs_ready;
  wire [3:0] constant472_outs;
  wire  constant472_outs_valid;
  wire  constant472_outs_ready;
  wire [4:0] extsi152_outs;
  wire  extsi152_outs_valid;
  wire  extsi152_outs_ready;
  wire [0:0] cmpi4_result;
  wire  cmpi4_result_valid;
  wire  cmpi4_result_ready;
  wire [0:0] fork15_outs_0;
  wire  fork15_outs_0_valid;
  wire  fork15_outs_0_ready;
  wire [0:0] fork15_outs_1;
  wire  fork15_outs_1_valid;
  wire  fork15_outs_1_ready;
  wire [0:0] fork15_outs_2;
  wire  fork15_outs_2_valid;
  wire  fork15_outs_2_ready;
  wire [0:0] fork15_outs_3;
  wire  fork15_outs_3_valid;
  wire  fork15_outs_3_ready;
  wire [0:0] fork15_outs_4;
  wire  fork15_outs_4_valid;
  wire  fork15_outs_4_ready;
  wire [0:0] fork15_outs_5;
  wire  fork15_outs_5_valid;
  wire  fork15_outs_5_ready;
  wire [0:0] fork15_outs_6;
  wire  fork15_outs_6_valid;
  wire  fork15_outs_6_ready;
  wire [0:0] fork15_outs_7;
  wire  fork15_outs_7_valid;
  wire  fork15_outs_7_ready;
  wire [0:0] fork15_outs_8;
  wire  fork15_outs_8_valid;
  wire  fork15_outs_8_ready;
  wire [35:0] cond_br68_trueOut;
  wire  cond_br68_trueOut_valid;
  wire  cond_br68_trueOut_ready;
  wire [35:0] cond_br68_falseOut;
  wire  cond_br68_falseOut_valid;
  wire  cond_br68_falseOut_ready;
  wire [36:0] extsi153_outs;
  wire  extsi153_outs_valid;
  wire  extsi153_outs_ready;
  wire [32:0] cond_br69_trueOut;
  wire  cond_br69_trueOut_valid;
  wire  cond_br69_trueOut_ready;
  wire [32:0] cond_br69_falseOut;
  wire  cond_br69_falseOut_valid;
  wire  cond_br69_falseOut_ready;
  wire [26:0] cond_br70_trueOut;
  wire  cond_br70_trueOut_valid;
  wire  cond_br70_trueOut_ready;
  wire [26:0] cond_br70_falseOut;
  wire  cond_br70_falseOut_valid;
  wire  cond_br70_falseOut_ready;
  wire [21:0] cond_br71_trueOut;
  wire  cond_br71_trueOut_valid;
  wire  cond_br71_trueOut_ready;
  wire [21:0] cond_br71_falseOut;
  wire  cond_br71_falseOut_valid;
  wire  cond_br71_falseOut_ready;
  wire [16:0] cond_br72_trueOut;
  wire  cond_br72_trueOut_valid;
  wire  cond_br72_trueOut_ready;
  wire [16:0] cond_br72_falseOut;
  wire  cond_br72_falseOut_valid;
  wire  cond_br72_falseOut_ready;
  wire [11:0] cond_br73_trueOut;
  wire  cond_br73_trueOut_valid;
  wire  cond_br73_trueOut_ready;
  wire [11:0] cond_br73_falseOut;
  wire  cond_br73_falseOut_valid;
  wire  cond_br73_falseOut_ready;
  wire [6:0] buffer18_outs;
  wire  buffer18_outs_valid;
  wire  buffer18_outs_ready;
  wire [6:0] buffer19_outs;
  wire  buffer19_outs_valid;
  wire  buffer19_outs_ready;
  wire [6:0] cond_br74_trueOut;
  wire  cond_br74_trueOut_valid;
  wire  cond_br74_trueOut_ready;
  wire [6:0] cond_br74_falseOut;
  wire  cond_br74_falseOut_valid;
  wire  cond_br74_falseOut_ready;
  wire  cond_br75_trueOut_valid;
  wire  cond_br75_trueOut_ready;
  wire  cond_br75_falseOut_valid;
  wire  cond_br75_falseOut_ready;
  wire [4:0] cond_br76_trueOut;
  wire  cond_br76_trueOut_valid;
  wire  cond_br76_trueOut_ready;
  wire [4:0] cond_br76_falseOut;
  wire  cond_br76_falseOut_valid;
  wire  cond_br76_falseOut_ready;
  wire [4:0] buffer26_outs;
  wire  buffer26_outs_valid;
  wire  buffer26_outs_ready;
  wire [4:0] buffer27_outs;
  wire  buffer27_outs_valid;
  wire  buffer27_outs_ready;
  wire [4:0] fork16_outs_0;
  wire  fork16_outs_0_valid;
  wire  fork16_outs_0_ready;
  wire [4:0] fork16_outs_1;
  wire  fork16_outs_1_valid;
  wire  fork16_outs_1_ready;
  wire  buffer28_outs_valid;
  wire  buffer28_outs_ready;
  wire  buffer29_outs_valid;
  wire  buffer29_outs_ready;
  wire  fork17_outs_0_valid;
  wire  fork17_outs_0_ready;
  wire  fork17_outs_1_valid;
  wire  fork17_outs_1_ready;
  wire  fork17_outs_2_valid;
  wire  fork17_outs_2_ready;
  wire  fork17_outs_3_valid;
  wire  fork17_outs_3_ready;
  wire  fork17_outs_4_valid;
  wire  fork17_outs_4_ready;
  wire  fork17_outs_5_valid;
  wire  fork17_outs_5_ready;
  wire  fork17_outs_6_valid;
  wire  fork17_outs_6_ready;
  wire [35:0] constant473_outs;
  wire  constant473_outs_valid;
  wire  constant473_outs_ready;
  wire [32:0] constant259_outs;
  wire  constant259_outs_valid;
  wire  constant259_outs_ready;
  wire [26:0] constant260_outs;
  wire  constant260_outs_valid;
  wire  constant260_outs_ready;
  wire [21:0] constant261_outs;
  wire  constant261_outs_valid;
  wire  constant261_outs_ready;
  wire [16:0] constant262_outs;
  wire  constant262_outs_valid;
  wire  constant262_outs_ready;
  wire [11:0] constant263_outs;
  wire  constant263_outs_valid;
  wire  constant263_outs_ready;
  wire  source6_outs_valid;
  wire  source6_outs_ready;
  wire [3:0] constant474_outs;
  wire  constant474_outs_valid;
  wire  constant474_outs_ready;
  wire [4:0] extsi154_outs;
  wire  extsi154_outs_valid;
  wire  extsi154_outs_ready;
  wire [0:0] cmpi5_result;
  wire  cmpi5_result_valid;
  wire  cmpi5_result_ready;
  wire [0:0] fork18_outs_0;
  wire  fork18_outs_0_valid;
  wire  fork18_outs_0_ready;
  wire [0:0] fork18_outs_1;
  wire  fork18_outs_1_valid;
  wire  fork18_outs_1_ready;
  wire [0:0] fork18_outs_2;
  wire  fork18_outs_2_valid;
  wire  fork18_outs_2_ready;
  wire [0:0] fork18_outs_3;
  wire  fork18_outs_3_valid;
  wire  fork18_outs_3_ready;
  wire [0:0] fork18_outs_4;
  wire  fork18_outs_4_valid;
  wire  fork18_outs_4_ready;
  wire [0:0] fork18_outs_5;
  wire  fork18_outs_5_valid;
  wire  fork18_outs_5_ready;
  wire [0:0] fork18_outs_6;
  wire  fork18_outs_6_valid;
  wire  fork18_outs_6_ready;
  wire [0:0] fork18_outs_7;
  wire  fork18_outs_7_valid;
  wire  fork18_outs_7_ready;
  wire [0:0] fork18_outs_8;
  wire  fork18_outs_8_valid;
  wire  fork18_outs_8_ready;
  wire [35:0] cond_br77_trueOut;
  wire  cond_br77_trueOut_valid;
  wire  cond_br77_trueOut_ready;
  wire [35:0] cond_br77_falseOut;
  wire  cond_br77_falseOut_valid;
  wire  cond_br77_falseOut_ready;
  wire [36:0] extsi155_outs;
  wire  extsi155_outs_valid;
  wire  extsi155_outs_ready;
  wire [32:0] cond_br78_trueOut;
  wire  cond_br78_trueOut_valid;
  wire  cond_br78_trueOut_ready;
  wire [32:0] cond_br78_falseOut;
  wire  cond_br78_falseOut_valid;
  wire  cond_br78_falseOut_ready;
  wire [26:0] cond_br79_trueOut;
  wire  cond_br79_trueOut_valid;
  wire  cond_br79_trueOut_ready;
  wire [26:0] cond_br79_falseOut;
  wire  cond_br79_falseOut_valid;
  wire  cond_br79_falseOut_ready;
  wire [21:0] cond_br80_trueOut;
  wire  cond_br80_trueOut_valid;
  wire  cond_br80_trueOut_ready;
  wire [21:0] cond_br80_falseOut;
  wire  cond_br80_falseOut_valid;
  wire  cond_br80_falseOut_ready;
  wire [16:0] cond_br81_trueOut;
  wire  cond_br81_trueOut_valid;
  wire  cond_br81_trueOut_ready;
  wire [16:0] cond_br81_falseOut;
  wire  cond_br81_falseOut_valid;
  wire  cond_br81_falseOut_ready;
  wire [11:0] cond_br82_trueOut;
  wire  cond_br82_trueOut_valid;
  wire  cond_br82_trueOut_ready;
  wire [11:0] cond_br82_falseOut;
  wire  cond_br82_falseOut_valid;
  wire  cond_br82_falseOut_ready;
  wire [6:0] buffer24_outs;
  wire  buffer24_outs_valid;
  wire  buffer24_outs_ready;
  wire [6:0] buffer25_outs;
  wire  buffer25_outs_valid;
  wire  buffer25_outs_ready;
  wire [6:0] cond_br83_trueOut;
  wire  cond_br83_trueOut_valid;
  wire  cond_br83_trueOut_ready;
  wire [6:0] cond_br83_falseOut;
  wire  cond_br83_falseOut_valid;
  wire  cond_br83_falseOut_ready;
  wire  cond_br84_trueOut_valid;
  wire  cond_br84_trueOut_ready;
  wire  cond_br84_falseOut_valid;
  wire  cond_br84_falseOut_ready;
  wire [4:0] cond_br85_trueOut;
  wire  cond_br85_trueOut_valid;
  wire  cond_br85_trueOut_ready;
  wire [4:0] cond_br85_falseOut;
  wire  cond_br85_falseOut_valid;
  wire  cond_br85_falseOut_ready;
  wire [4:0] buffer32_outs;
  wire  buffer32_outs_valid;
  wire  buffer32_outs_ready;
  wire [4:0] buffer33_outs;
  wire  buffer33_outs_valid;
  wire  buffer33_outs_ready;
  wire [4:0] fork19_outs_0;
  wire  fork19_outs_0_valid;
  wire  fork19_outs_0_ready;
  wire [4:0] fork19_outs_1;
  wire  fork19_outs_1_valid;
  wire  fork19_outs_1_ready;
  wire  buffer34_outs_valid;
  wire  buffer34_outs_ready;
  wire  buffer35_outs_valid;
  wire  buffer35_outs_ready;
  wire  fork20_outs_0_valid;
  wire  fork20_outs_0_ready;
  wire  fork20_outs_1_valid;
  wire  fork20_outs_1_ready;
  wire  fork20_outs_2_valid;
  wire  fork20_outs_2_ready;
  wire  fork20_outs_3_valid;
  wire  fork20_outs_3_ready;
  wire  fork20_outs_4_valid;
  wire  fork20_outs_4_ready;
  wire  fork20_outs_5_valid;
  wire  fork20_outs_5_ready;
  wire  fork20_outs_6_valid;
  wire  fork20_outs_6_ready;
  wire [35:0] constant475_outs;
  wire  constant475_outs_valid;
  wire  constant475_outs_ready;
  wire [31:0] constant476_outs;
  wire  constant476_outs_valid;
  wire  constant476_outs_ready;
  wire [26:0] constant267_outs;
  wire  constant267_outs_valid;
  wire  constant267_outs_ready;
  wire [21:0] constant268_outs;
  wire  constant268_outs_valid;
  wire  constant268_outs_ready;
  wire [16:0] constant269_outs;
  wire  constant269_outs_valid;
  wire  constant269_outs_ready;
  wire [11:0] constant270_outs;
  wire  constant270_outs_valid;
  wire  constant270_outs_ready;
  wire  source7_outs_valid;
  wire  source7_outs_ready;
  wire [3:0] constant477_outs;
  wire  constant477_outs_valid;
  wire  constant477_outs_ready;
  wire [4:0] extsi156_outs;
  wire  extsi156_outs_valid;
  wire  extsi156_outs_ready;
  wire [0:0] cmpi6_result;
  wire  cmpi6_result_valid;
  wire  cmpi6_result_ready;
  wire [0:0] fork21_outs_0;
  wire  fork21_outs_0_valid;
  wire  fork21_outs_0_ready;
  wire [0:0] fork21_outs_1;
  wire  fork21_outs_1_valid;
  wire  fork21_outs_1_ready;
  wire [0:0] fork21_outs_2;
  wire  fork21_outs_2_valid;
  wire  fork21_outs_2_ready;
  wire [0:0] fork21_outs_3;
  wire  fork21_outs_3_valid;
  wire  fork21_outs_3_ready;
  wire [0:0] fork21_outs_4;
  wire  fork21_outs_4_valid;
  wire  fork21_outs_4_ready;
  wire [0:0] fork21_outs_5;
  wire  fork21_outs_5_valid;
  wire  fork21_outs_5_ready;
  wire [0:0] fork21_outs_6;
  wire  fork21_outs_6_valid;
  wire  fork21_outs_6_ready;
  wire [0:0] fork21_outs_7;
  wire  fork21_outs_7_valid;
  wire  fork21_outs_7_ready;
  wire [0:0] fork21_outs_8;
  wire  fork21_outs_8_valid;
  wire  fork21_outs_8_ready;
  wire [35:0] cond_br86_trueOut;
  wire  cond_br86_trueOut_valid;
  wire  cond_br86_trueOut_ready;
  wire [35:0] cond_br86_falseOut;
  wire  cond_br86_falseOut_valid;
  wire  cond_br86_falseOut_ready;
  wire [36:0] extsi157_outs;
  wire  extsi157_outs_valid;
  wire  extsi157_outs_ready;
  wire [31:0] cond_br87_trueOut;
  wire  cond_br87_trueOut_valid;
  wire  cond_br87_trueOut_ready;
  wire [31:0] cond_br87_falseOut;
  wire  cond_br87_falseOut_valid;
  wire  cond_br87_falseOut_ready;
  wire [32:0] extsi158_outs;
  wire  extsi158_outs_valid;
  wire  extsi158_outs_ready;
  wire [26:0] cond_br88_trueOut;
  wire  cond_br88_trueOut_valid;
  wire  cond_br88_trueOut_ready;
  wire [26:0] cond_br88_falseOut;
  wire  cond_br88_falseOut_valid;
  wire  cond_br88_falseOut_ready;
  wire [21:0] cond_br89_trueOut;
  wire  cond_br89_trueOut_valid;
  wire  cond_br89_trueOut_ready;
  wire [21:0] cond_br89_falseOut;
  wire  cond_br89_falseOut_valid;
  wire  cond_br89_falseOut_ready;
  wire [16:0] cond_br90_trueOut;
  wire  cond_br90_trueOut_valid;
  wire  cond_br90_trueOut_ready;
  wire [16:0] cond_br90_falseOut;
  wire  cond_br90_falseOut_valid;
  wire  cond_br90_falseOut_ready;
  wire [11:0] cond_br91_trueOut;
  wire  cond_br91_trueOut_valid;
  wire  cond_br91_trueOut_ready;
  wire [11:0] cond_br91_falseOut;
  wire  cond_br91_falseOut_valid;
  wire  cond_br91_falseOut_ready;
  wire [6:0] buffer30_outs;
  wire  buffer30_outs_valid;
  wire  buffer30_outs_ready;
  wire [6:0] buffer31_outs;
  wire  buffer31_outs_valid;
  wire  buffer31_outs_ready;
  wire [6:0] cond_br92_trueOut;
  wire  cond_br92_trueOut_valid;
  wire  cond_br92_trueOut_ready;
  wire [6:0] cond_br92_falseOut;
  wire  cond_br92_falseOut_valid;
  wire  cond_br92_falseOut_ready;
  wire  cond_br93_trueOut_valid;
  wire  cond_br93_trueOut_ready;
  wire  cond_br93_falseOut_valid;
  wire  cond_br93_falseOut_ready;
  wire [4:0] cond_br94_trueOut;
  wire  cond_br94_trueOut_valid;
  wire  cond_br94_trueOut_ready;
  wire [4:0] cond_br94_falseOut;
  wire  cond_br94_falseOut_valid;
  wire  cond_br94_falseOut_ready;
  wire [4:0] buffer38_outs;
  wire  buffer38_outs_valid;
  wire  buffer38_outs_ready;
  wire [4:0] buffer39_outs;
  wire  buffer39_outs_valid;
  wire  buffer39_outs_ready;
  wire [4:0] fork22_outs_0;
  wire  fork22_outs_0_valid;
  wire  fork22_outs_0_ready;
  wire [4:0] fork22_outs_1;
  wire  fork22_outs_1_valid;
  wire  fork22_outs_1_ready;
  wire  buffer40_outs_valid;
  wire  buffer40_outs_ready;
  wire  buffer41_outs_valid;
  wire  buffer41_outs_ready;
  wire  fork23_outs_0_valid;
  wire  fork23_outs_0_ready;
  wire  fork23_outs_1_valid;
  wire  fork23_outs_1_ready;
  wire  fork23_outs_2_valid;
  wire  fork23_outs_2_ready;
  wire  fork23_outs_3_valid;
  wire  fork23_outs_3_ready;
  wire  fork23_outs_4_valid;
  wire  fork23_outs_4_ready;
  wire  fork23_outs_5_valid;
  wire  fork23_outs_5_ready;
  wire  fork23_outs_6_valid;
  wire  fork23_outs_6_ready;
  wire [36:0] constant272_outs;
  wire  constant272_outs_valid;
  wire  constant272_outs_ready;
  wire [31:0] constant478_outs;
  wire  constant478_outs_valid;
  wire  constant478_outs_ready;
  wire [26:0] constant274_outs;
  wire  constant274_outs_valid;
  wire  constant274_outs_ready;
  wire [18:0] constant479_outs;
  wire  constant479_outs_valid;
  wire  constant479_outs_ready;
  wire [16:0] constant276_outs;
  wire  constant276_outs_valid;
  wire  constant276_outs_ready;
  wire [11:0] constant277_outs;
  wire  constant277_outs_valid;
  wire  constant277_outs_ready;
  wire  source8_outs_valid;
  wire  source8_outs_ready;
  wire [3:0] constant480_outs;
  wire  constant480_outs_valid;
  wire  constant480_outs_ready;
  wire [4:0] extsi159_outs;
  wire  extsi159_outs_valid;
  wire  extsi159_outs_ready;
  wire [0:0] cmpi7_result;
  wire  cmpi7_result_valid;
  wire  cmpi7_result_ready;
  wire [0:0] fork24_outs_0;
  wire  fork24_outs_0_valid;
  wire  fork24_outs_0_ready;
  wire [0:0] fork24_outs_1;
  wire  fork24_outs_1_valid;
  wire  fork24_outs_1_ready;
  wire [0:0] fork24_outs_2;
  wire  fork24_outs_2_valid;
  wire  fork24_outs_2_ready;
  wire [0:0] fork24_outs_3;
  wire  fork24_outs_3_valid;
  wire  fork24_outs_3_ready;
  wire [0:0] fork24_outs_4;
  wire  fork24_outs_4_valid;
  wire  fork24_outs_4_ready;
  wire [0:0] fork24_outs_5;
  wire  fork24_outs_5_valid;
  wire  fork24_outs_5_ready;
  wire [0:0] fork24_outs_6;
  wire  fork24_outs_6_valid;
  wire  fork24_outs_6_ready;
  wire [0:0] fork24_outs_7;
  wire  fork24_outs_7_valid;
  wire  fork24_outs_7_ready;
  wire [0:0] fork24_outs_8;
  wire  fork24_outs_8_valid;
  wire  fork24_outs_8_ready;
  wire [36:0] cond_br95_trueOut;
  wire  cond_br95_trueOut_valid;
  wire  cond_br95_trueOut_ready;
  wire [36:0] cond_br95_falseOut;
  wire  cond_br95_falseOut_valid;
  wire  cond_br95_falseOut_ready;
  wire [31:0] cond_br96_trueOut;
  wire  cond_br96_trueOut_valid;
  wire  cond_br96_trueOut_ready;
  wire [31:0] cond_br96_falseOut;
  wire  cond_br96_falseOut_valid;
  wire  cond_br96_falseOut_ready;
  wire [32:0] extsi160_outs;
  wire  extsi160_outs_valid;
  wire  extsi160_outs_ready;
  wire [26:0] cond_br97_trueOut;
  wire  cond_br97_trueOut_valid;
  wire  cond_br97_trueOut_ready;
  wire [26:0] cond_br97_falseOut;
  wire  cond_br97_falseOut_valid;
  wire  cond_br97_falseOut_ready;
  wire [18:0] cond_br98_trueOut;
  wire  cond_br98_trueOut_valid;
  wire  cond_br98_trueOut_ready;
  wire [18:0] cond_br98_falseOut;
  wire  cond_br98_falseOut_valid;
  wire  cond_br98_falseOut_ready;
  wire [21:0] extsi161_outs;
  wire  extsi161_outs_valid;
  wire  extsi161_outs_ready;
  wire [16:0] cond_br99_trueOut;
  wire  cond_br99_trueOut_valid;
  wire  cond_br99_trueOut_ready;
  wire [16:0] cond_br99_falseOut;
  wire  cond_br99_falseOut_valid;
  wire  cond_br99_falseOut_ready;
  wire [11:0] cond_br100_trueOut;
  wire  cond_br100_trueOut_valid;
  wire  cond_br100_trueOut_ready;
  wire [11:0] cond_br100_falseOut;
  wire  cond_br100_falseOut_valid;
  wire  cond_br100_falseOut_ready;
  wire [6:0] buffer36_outs;
  wire  buffer36_outs_valid;
  wire  buffer36_outs_ready;
  wire [6:0] buffer37_outs;
  wire  buffer37_outs_valid;
  wire  buffer37_outs_ready;
  wire [6:0] cond_br101_trueOut;
  wire  cond_br101_trueOut_valid;
  wire  cond_br101_trueOut_ready;
  wire [6:0] cond_br101_falseOut;
  wire  cond_br101_falseOut_valid;
  wire  cond_br101_falseOut_ready;
  wire  cond_br102_trueOut_valid;
  wire  cond_br102_trueOut_ready;
  wire  cond_br102_falseOut_valid;
  wire  cond_br102_falseOut_ready;
  wire [4:0] cond_br103_trueOut;
  wire  cond_br103_trueOut_valid;
  wire  cond_br103_trueOut_ready;
  wire [4:0] cond_br103_falseOut;
  wire  cond_br103_falseOut_valid;
  wire  cond_br103_falseOut_ready;
  wire [4:0] buffer44_outs;
  wire  buffer44_outs_valid;
  wire  buffer44_outs_ready;
  wire [4:0] buffer45_outs;
  wire  buffer45_outs_valid;
  wire  buffer45_outs_ready;
  wire [4:0] fork25_outs_0;
  wire  fork25_outs_0_valid;
  wire  fork25_outs_0_ready;
  wire [4:0] fork25_outs_1;
  wire  fork25_outs_1_valid;
  wire  fork25_outs_1_ready;
  wire  buffer46_outs_valid;
  wire  buffer46_outs_ready;
  wire  buffer47_outs_valid;
  wire  buffer47_outs_ready;
  wire  fork26_outs_0_valid;
  wire  fork26_outs_0_ready;
  wire  fork26_outs_1_valid;
  wire  fork26_outs_1_ready;
  wire  fork26_outs_2_valid;
  wire  fork26_outs_2_ready;
  wire  fork26_outs_3_valid;
  wire  fork26_outs_3_ready;
  wire  fork26_outs_4_valid;
  wire  fork26_outs_4_ready;
  wire  fork26_outs_5_valid;
  wire  fork26_outs_5_ready;
  wire  fork26_outs_6_valid;
  wire  fork26_outs_6_ready;
  wire [36:0] constant279_outs;
  wire  constant279_outs_valid;
  wire  constant279_outs_ready;
  wire [31:0] constant481_outs;
  wire  constant481_outs_valid;
  wire  constant481_outs_ready;
  wire [26:0] constant281_outs;
  wire  constant281_outs_valid;
  wire  constant281_outs_ready;
  wire [19:0] constant482_outs;
  wire  constant482_outs_valid;
  wire  constant482_outs_ready;
  wire [15:0] constant483_outs;
  wire  constant483_outs_valid;
  wire  constant483_outs_ready;
  wire [11:0] constant284_outs;
  wire  constant284_outs_valid;
  wire  constant284_outs_ready;
  wire  source9_outs_valid;
  wire  source9_outs_ready;
  wire [4:0] constant484_outs;
  wire  constant484_outs_valid;
  wire  constant484_outs_ready;
  wire [0:0] cmpi8_result;
  wire  cmpi8_result_valid;
  wire  cmpi8_result_ready;
  wire [0:0] fork27_outs_0;
  wire  fork27_outs_0_valid;
  wire  fork27_outs_0_ready;
  wire [0:0] fork27_outs_1;
  wire  fork27_outs_1_valid;
  wire  fork27_outs_1_ready;
  wire [0:0] fork27_outs_2;
  wire  fork27_outs_2_valid;
  wire  fork27_outs_2_ready;
  wire [0:0] fork27_outs_3;
  wire  fork27_outs_3_valid;
  wire  fork27_outs_3_ready;
  wire [0:0] fork27_outs_4;
  wire  fork27_outs_4_valid;
  wire  fork27_outs_4_ready;
  wire [0:0] fork27_outs_5;
  wire  fork27_outs_5_valid;
  wire  fork27_outs_5_ready;
  wire [0:0] fork27_outs_6;
  wire  fork27_outs_6_valid;
  wire  fork27_outs_6_ready;
  wire [0:0] fork27_outs_7;
  wire  fork27_outs_7_valid;
  wire  fork27_outs_7_ready;
  wire [0:0] fork27_outs_8;
  wire  fork27_outs_8_valid;
  wire  fork27_outs_8_ready;
  wire [36:0] cond_br104_trueOut;
  wire  cond_br104_trueOut_valid;
  wire  cond_br104_trueOut_ready;
  wire [36:0] cond_br104_falseOut;
  wire  cond_br104_falseOut_valid;
  wire  cond_br104_falseOut_ready;
  wire [31:0] cond_br105_trueOut;
  wire  cond_br105_trueOut_valid;
  wire  cond_br105_trueOut_ready;
  wire [31:0] cond_br105_falseOut;
  wire  cond_br105_falseOut_valid;
  wire  cond_br105_falseOut_ready;
  wire [32:0] extsi162_outs;
  wire  extsi162_outs_valid;
  wire  extsi162_outs_ready;
  wire [26:0] cond_br106_trueOut;
  wire  cond_br106_trueOut_valid;
  wire  cond_br106_trueOut_ready;
  wire [26:0] cond_br106_falseOut;
  wire  cond_br106_falseOut_valid;
  wire  cond_br106_falseOut_ready;
  wire [19:0] cond_br107_trueOut;
  wire  cond_br107_trueOut_valid;
  wire  cond_br107_trueOut_ready;
  wire [19:0] cond_br107_falseOut;
  wire  cond_br107_falseOut_valid;
  wire  cond_br107_falseOut_ready;
  wire [21:0] extsi163_outs;
  wire  extsi163_outs_valid;
  wire  extsi163_outs_ready;
  wire [15:0] cond_br108_trueOut;
  wire  cond_br108_trueOut_valid;
  wire  cond_br108_trueOut_ready;
  wire [15:0] cond_br108_falseOut;
  wire  cond_br108_falseOut_valid;
  wire  cond_br108_falseOut_ready;
  wire [16:0] extsi164_outs;
  wire  extsi164_outs_valid;
  wire  extsi164_outs_ready;
  wire [11:0] cond_br109_trueOut;
  wire  cond_br109_trueOut_valid;
  wire  cond_br109_trueOut_ready;
  wire [11:0] cond_br109_falseOut;
  wire  cond_br109_falseOut_valid;
  wire  cond_br109_falseOut_ready;
  wire [6:0] buffer42_outs;
  wire  buffer42_outs_valid;
  wire  buffer42_outs_ready;
  wire [6:0] buffer43_outs;
  wire  buffer43_outs_valid;
  wire  buffer43_outs_ready;
  wire [6:0] cond_br110_trueOut;
  wire  cond_br110_trueOut_valid;
  wire  cond_br110_trueOut_ready;
  wire [6:0] cond_br110_falseOut;
  wire  cond_br110_falseOut_valid;
  wire  cond_br110_falseOut_ready;
  wire  cond_br111_trueOut_valid;
  wire  cond_br111_trueOut_ready;
  wire  cond_br111_falseOut_valid;
  wire  cond_br111_falseOut_ready;
  wire [4:0] cond_br112_trueOut;
  wire  cond_br112_trueOut_valid;
  wire  cond_br112_trueOut_ready;
  wire [4:0] cond_br112_falseOut;
  wire  cond_br112_falseOut_valid;
  wire  cond_br112_falseOut_ready;
  wire [4:0] buffer50_outs;
  wire  buffer50_outs_valid;
  wire  buffer50_outs_ready;
  wire [4:0] buffer51_outs;
  wire  buffer51_outs_valid;
  wire  buffer51_outs_ready;
  wire [4:0] fork28_outs_0;
  wire  fork28_outs_0_valid;
  wire  fork28_outs_0_ready;
  wire [4:0] fork28_outs_1;
  wire  fork28_outs_1_valid;
  wire  fork28_outs_1_ready;
  wire  buffer52_outs_valid;
  wire  buffer52_outs_ready;
  wire  buffer53_outs_valid;
  wire  buffer53_outs_ready;
  wire  fork29_outs_0_valid;
  wire  fork29_outs_0_ready;
  wire  fork29_outs_1_valid;
  wire  fork29_outs_1_ready;
  wire  fork29_outs_2_valid;
  wire  fork29_outs_2_ready;
  wire  fork29_outs_3_valid;
  wire  fork29_outs_3_ready;
  wire  fork29_outs_4_valid;
  wire  fork29_outs_4_ready;
  wire  fork29_outs_5_valid;
  wire  fork29_outs_5_ready;
  wire  fork29_outs_6_valid;
  wire  fork29_outs_6_ready;
  wire [36:0] constant286_outs;
  wire  constant286_outs_valid;
  wire  constant286_outs_ready;
  wire [31:0] constant485_outs;
  wire  constant485_outs_valid;
  wire  constant485_outs_ready;
  wire [26:0] constant288_outs;
  wire  constant288_outs_valid;
  wire  constant288_outs_ready;
  wire [20:0] constant486_outs;
  wire  constant486_outs_valid;
  wire  constant486_outs_ready;
  wire [15:0] constant487_outs;
  wire  constant487_outs_valid;
  wire  constant487_outs_ready;
  wire [11:0] constant291_outs;
  wire  constant291_outs_valid;
  wire  constant291_outs_ready;
  wire  source10_outs_valid;
  wire  source10_outs_ready;
  wire [4:0] constant488_outs;
  wire  constant488_outs_valid;
  wire  constant488_outs_ready;
  wire [0:0] cmpi9_result;
  wire  cmpi9_result_valid;
  wire  cmpi9_result_ready;
  wire [0:0] fork30_outs_0;
  wire  fork30_outs_0_valid;
  wire  fork30_outs_0_ready;
  wire [0:0] fork30_outs_1;
  wire  fork30_outs_1_valid;
  wire  fork30_outs_1_ready;
  wire [0:0] fork30_outs_2;
  wire  fork30_outs_2_valid;
  wire  fork30_outs_2_ready;
  wire [0:0] fork30_outs_3;
  wire  fork30_outs_3_valid;
  wire  fork30_outs_3_ready;
  wire [0:0] fork30_outs_4;
  wire  fork30_outs_4_valid;
  wire  fork30_outs_4_ready;
  wire [0:0] fork30_outs_5;
  wire  fork30_outs_5_valid;
  wire  fork30_outs_5_ready;
  wire [0:0] fork30_outs_6;
  wire  fork30_outs_6_valid;
  wire  fork30_outs_6_ready;
  wire [0:0] fork30_outs_7;
  wire  fork30_outs_7_valid;
  wire  fork30_outs_7_ready;
  wire [0:0] fork30_outs_8;
  wire  fork30_outs_8_valid;
  wire  fork30_outs_8_ready;
  wire [36:0] cond_br113_trueOut;
  wire  cond_br113_trueOut_valid;
  wire  cond_br113_trueOut_ready;
  wire [36:0] cond_br113_falseOut;
  wire  cond_br113_falseOut_valid;
  wire  cond_br113_falseOut_ready;
  wire [31:0] cond_br114_trueOut;
  wire  cond_br114_trueOut_valid;
  wire  cond_br114_trueOut_ready;
  wire [31:0] cond_br114_falseOut;
  wire  cond_br114_falseOut_valid;
  wire  cond_br114_falseOut_ready;
  wire [32:0] extsi165_outs;
  wire  extsi165_outs_valid;
  wire  extsi165_outs_ready;
  wire [26:0] cond_br115_trueOut;
  wire  cond_br115_trueOut_valid;
  wire  cond_br115_trueOut_ready;
  wire [26:0] cond_br115_falseOut;
  wire  cond_br115_falseOut_valid;
  wire  cond_br115_falseOut_ready;
  wire [20:0] cond_br116_trueOut;
  wire  cond_br116_trueOut_valid;
  wire  cond_br116_trueOut_ready;
  wire [20:0] cond_br116_falseOut;
  wire  cond_br116_falseOut_valid;
  wire  cond_br116_falseOut_ready;
  wire [21:0] extsi166_outs;
  wire  extsi166_outs_valid;
  wire  extsi166_outs_ready;
  wire [15:0] cond_br117_trueOut;
  wire  cond_br117_trueOut_valid;
  wire  cond_br117_trueOut_ready;
  wire [15:0] cond_br117_falseOut;
  wire  cond_br117_falseOut_valid;
  wire  cond_br117_falseOut_ready;
  wire [16:0] extsi167_outs;
  wire  extsi167_outs_valid;
  wire  extsi167_outs_ready;
  wire [11:0] cond_br118_trueOut;
  wire  cond_br118_trueOut_valid;
  wire  cond_br118_trueOut_ready;
  wire [11:0] cond_br118_falseOut;
  wire  cond_br118_falseOut_valid;
  wire  cond_br118_falseOut_ready;
  wire [6:0] buffer48_outs;
  wire  buffer48_outs_valid;
  wire  buffer48_outs_ready;
  wire [6:0] buffer49_outs;
  wire  buffer49_outs_valid;
  wire  buffer49_outs_ready;
  wire [6:0] cond_br119_trueOut;
  wire  cond_br119_trueOut_valid;
  wire  cond_br119_trueOut_ready;
  wire [6:0] cond_br119_falseOut;
  wire  cond_br119_falseOut_valid;
  wire  cond_br119_falseOut_ready;
  wire  cond_br120_trueOut_valid;
  wire  cond_br120_trueOut_ready;
  wire  cond_br120_falseOut_valid;
  wire  cond_br120_falseOut_ready;
  wire [4:0] cond_br121_trueOut;
  wire  cond_br121_trueOut_valid;
  wire  cond_br121_trueOut_ready;
  wire [4:0] cond_br121_falseOut;
  wire  cond_br121_falseOut_valid;
  wire  cond_br121_falseOut_ready;
  wire [4:0] buffer56_outs;
  wire  buffer56_outs_valid;
  wire  buffer56_outs_ready;
  wire [4:0] buffer57_outs;
  wire  buffer57_outs_valid;
  wire  buffer57_outs_ready;
  wire [4:0] fork31_outs_0;
  wire  fork31_outs_0_valid;
  wire  fork31_outs_0_ready;
  wire [4:0] fork31_outs_1;
  wire  fork31_outs_1_valid;
  wire  fork31_outs_1_ready;
  wire  buffer58_outs_valid;
  wire  buffer58_outs_ready;
  wire  buffer59_outs_valid;
  wire  buffer59_outs_ready;
  wire  fork32_outs_0_valid;
  wire  fork32_outs_0_ready;
  wire  fork32_outs_1_valid;
  wire  fork32_outs_1_ready;
  wire  fork32_outs_2_valid;
  wire  fork32_outs_2_ready;
  wire  fork32_outs_3_valid;
  wire  fork32_outs_3_ready;
  wire  fork32_outs_4_valid;
  wire  fork32_outs_4_ready;
  wire  fork32_outs_5_valid;
  wire  fork32_outs_5_ready;
  wire  fork32_outs_6_valid;
  wire  fork32_outs_6_ready;
  wire [36:0] constant293_outs;
  wire  constant293_outs_valid;
  wire  constant293_outs_ready;
  wire [31:0] constant489_outs;
  wire  constant489_outs_valid;
  wire  constant489_outs_ready;
  wire [26:0] constant295_outs;
  wire  constant295_outs_valid;
  wire  constant295_outs_ready;
  wire [20:0] constant490_outs;
  wire  constant490_outs_valid;
  wire  constant490_outs_ready;
  wire [14:0] constant491_outs;
  wire  constant491_outs_valid;
  wire  constant491_outs_ready;
  wire [11:0] constant298_outs;
  wire  constant298_outs_valid;
  wire  constant298_outs_ready;
  wire  source11_outs_valid;
  wire  source11_outs_ready;
  wire [4:0] constant492_outs;
  wire  constant492_outs_valid;
  wire  constant492_outs_ready;
  wire [0:0] cmpi10_result;
  wire  cmpi10_result_valid;
  wire  cmpi10_result_ready;
  wire [0:0] fork33_outs_0;
  wire  fork33_outs_0_valid;
  wire  fork33_outs_0_ready;
  wire [0:0] fork33_outs_1;
  wire  fork33_outs_1_valid;
  wire  fork33_outs_1_ready;
  wire [0:0] fork33_outs_2;
  wire  fork33_outs_2_valid;
  wire  fork33_outs_2_ready;
  wire [0:0] fork33_outs_3;
  wire  fork33_outs_3_valid;
  wire  fork33_outs_3_ready;
  wire [0:0] fork33_outs_4;
  wire  fork33_outs_4_valid;
  wire  fork33_outs_4_ready;
  wire [0:0] fork33_outs_5;
  wire  fork33_outs_5_valid;
  wire  fork33_outs_5_ready;
  wire [0:0] fork33_outs_6;
  wire  fork33_outs_6_valid;
  wire  fork33_outs_6_ready;
  wire [0:0] fork33_outs_7;
  wire  fork33_outs_7_valid;
  wire  fork33_outs_7_ready;
  wire [0:0] fork33_outs_8;
  wire  fork33_outs_8_valid;
  wire  fork33_outs_8_ready;
  wire [36:0] cond_br122_trueOut;
  wire  cond_br122_trueOut_valid;
  wire  cond_br122_trueOut_ready;
  wire [36:0] cond_br122_falseOut;
  wire  cond_br122_falseOut_valid;
  wire  cond_br122_falseOut_ready;
  wire [31:0] cond_br123_trueOut;
  wire  cond_br123_trueOut_valid;
  wire  cond_br123_trueOut_ready;
  wire [31:0] cond_br123_falseOut;
  wire  cond_br123_falseOut_valid;
  wire  cond_br123_falseOut_ready;
  wire [32:0] extsi168_outs;
  wire  extsi168_outs_valid;
  wire  extsi168_outs_ready;
  wire [26:0] cond_br124_trueOut;
  wire  cond_br124_trueOut_valid;
  wire  cond_br124_trueOut_ready;
  wire [26:0] cond_br124_falseOut;
  wire  cond_br124_falseOut_valid;
  wire  cond_br124_falseOut_ready;
  wire [20:0] cond_br125_trueOut;
  wire  cond_br125_trueOut_valid;
  wire  cond_br125_trueOut_ready;
  wire [20:0] cond_br125_falseOut;
  wire  cond_br125_falseOut_valid;
  wire  cond_br125_falseOut_ready;
  wire [21:0] extsi169_outs;
  wire  extsi169_outs_valid;
  wire  extsi169_outs_ready;
  wire [14:0] cond_br126_trueOut;
  wire  cond_br126_trueOut_valid;
  wire  cond_br126_trueOut_ready;
  wire [14:0] cond_br126_falseOut;
  wire  cond_br126_falseOut_valid;
  wire  cond_br126_falseOut_ready;
  wire [16:0] extsi170_outs;
  wire  extsi170_outs_valid;
  wire  extsi170_outs_ready;
  wire [11:0] cond_br127_trueOut;
  wire  cond_br127_trueOut_valid;
  wire  cond_br127_trueOut_ready;
  wire [11:0] cond_br127_falseOut;
  wire  cond_br127_falseOut_valid;
  wire  cond_br127_falseOut_ready;
  wire [6:0] buffer54_outs;
  wire  buffer54_outs_valid;
  wire  buffer54_outs_ready;
  wire [6:0] buffer55_outs;
  wire  buffer55_outs_valid;
  wire  buffer55_outs_ready;
  wire [6:0] cond_br128_trueOut;
  wire  cond_br128_trueOut_valid;
  wire  cond_br128_trueOut_ready;
  wire [6:0] cond_br128_falseOut;
  wire  cond_br128_falseOut_valid;
  wire  cond_br128_falseOut_ready;
  wire  cond_br129_trueOut_valid;
  wire  cond_br129_trueOut_ready;
  wire  cond_br129_falseOut_valid;
  wire  cond_br129_falseOut_ready;
  wire [4:0] cond_br130_trueOut;
  wire  cond_br130_trueOut_valid;
  wire  cond_br130_trueOut_ready;
  wire [4:0] cond_br130_falseOut;
  wire  cond_br130_falseOut_valid;
  wire  cond_br130_falseOut_ready;
  wire [4:0] buffer62_outs;
  wire  buffer62_outs_valid;
  wire  buffer62_outs_ready;
  wire [4:0] buffer63_outs;
  wire  buffer63_outs_valid;
  wire  buffer63_outs_ready;
  wire [4:0] fork34_outs_0;
  wire  fork34_outs_0_valid;
  wire  fork34_outs_0_ready;
  wire [4:0] fork34_outs_1;
  wire  fork34_outs_1_valid;
  wire  fork34_outs_1_ready;
  wire  buffer64_outs_valid;
  wire  buffer64_outs_ready;
  wire  buffer65_outs_valid;
  wire  buffer65_outs_ready;
  wire  fork35_outs_0_valid;
  wire  fork35_outs_0_ready;
  wire  fork35_outs_1_valid;
  wire  fork35_outs_1_ready;
  wire  fork35_outs_2_valid;
  wire  fork35_outs_2_ready;
  wire  fork35_outs_3_valid;
  wire  fork35_outs_3_ready;
  wire  fork35_outs_4_valid;
  wire  fork35_outs_4_ready;
  wire  fork35_outs_5_valid;
  wire  fork35_outs_5_ready;
  wire  fork35_outs_6_valid;
  wire  fork35_outs_6_ready;
  wire [36:0] constant300_outs;
  wire  constant300_outs_valid;
  wire  constant300_outs_ready;
  wire [30:0] constant493_outs;
  wire  constant493_outs_valid;
  wire  constant493_outs_ready;
  wire [26:0] constant302_outs;
  wire  constant302_outs_valid;
  wire  constant302_outs_ready;
  wire [20:0] constant494_outs;
  wire  constant494_outs_valid;
  wire  constant494_outs_ready;
  wire [12:0] constant495_outs;
  wire  constant495_outs_valid;
  wire  constant495_outs_ready;
  wire [11:0] constant305_outs;
  wire  constant305_outs_valid;
  wire  constant305_outs_ready;
  wire  source12_outs_valid;
  wire  source12_outs_ready;
  wire [4:0] constant496_outs;
  wire  constant496_outs_valid;
  wire  constant496_outs_ready;
  wire [0:0] cmpi11_result;
  wire  cmpi11_result_valid;
  wire  cmpi11_result_ready;
  wire [0:0] fork36_outs_0;
  wire  fork36_outs_0_valid;
  wire  fork36_outs_0_ready;
  wire [0:0] fork36_outs_1;
  wire  fork36_outs_1_valid;
  wire  fork36_outs_1_ready;
  wire [0:0] fork36_outs_2;
  wire  fork36_outs_2_valid;
  wire  fork36_outs_2_ready;
  wire [0:0] fork36_outs_3;
  wire  fork36_outs_3_valid;
  wire  fork36_outs_3_ready;
  wire [0:0] fork36_outs_4;
  wire  fork36_outs_4_valid;
  wire  fork36_outs_4_ready;
  wire [0:0] fork36_outs_5;
  wire  fork36_outs_5_valid;
  wire  fork36_outs_5_ready;
  wire [0:0] fork36_outs_6;
  wire  fork36_outs_6_valid;
  wire  fork36_outs_6_ready;
  wire [0:0] fork36_outs_7;
  wire  fork36_outs_7_valid;
  wire  fork36_outs_7_ready;
  wire [0:0] fork36_outs_8;
  wire  fork36_outs_8_valid;
  wire  fork36_outs_8_ready;
  wire [36:0] cond_br131_trueOut;
  wire  cond_br131_trueOut_valid;
  wire  cond_br131_trueOut_ready;
  wire [36:0] cond_br131_falseOut;
  wire  cond_br131_falseOut_valid;
  wire  cond_br131_falseOut_ready;
  wire [30:0] cond_br132_trueOut;
  wire  cond_br132_trueOut_valid;
  wire  cond_br132_trueOut_ready;
  wire [30:0] cond_br132_falseOut;
  wire  cond_br132_falseOut_valid;
  wire  cond_br132_falseOut_ready;
  wire [32:0] extsi171_outs;
  wire  extsi171_outs_valid;
  wire  extsi171_outs_ready;
  wire [26:0] cond_br133_trueOut;
  wire  cond_br133_trueOut_valid;
  wire  cond_br133_trueOut_ready;
  wire [26:0] cond_br133_falseOut;
  wire  cond_br133_falseOut_valid;
  wire  cond_br133_falseOut_ready;
  wire [20:0] cond_br134_trueOut;
  wire  cond_br134_trueOut_valid;
  wire  cond_br134_trueOut_ready;
  wire [20:0] cond_br134_falseOut;
  wire  cond_br134_falseOut_valid;
  wire  cond_br134_falseOut_ready;
  wire [21:0] extsi172_outs;
  wire  extsi172_outs_valid;
  wire  extsi172_outs_ready;
  wire [12:0] cond_br135_trueOut;
  wire  cond_br135_trueOut_valid;
  wire  cond_br135_trueOut_ready;
  wire [12:0] cond_br135_falseOut;
  wire  cond_br135_falseOut_valid;
  wire  cond_br135_falseOut_ready;
  wire [16:0] extsi173_outs;
  wire  extsi173_outs_valid;
  wire  extsi173_outs_ready;
  wire [11:0] cond_br136_trueOut;
  wire  cond_br136_trueOut_valid;
  wire  cond_br136_trueOut_ready;
  wire [11:0] cond_br136_falseOut;
  wire  cond_br136_falseOut_valid;
  wire  cond_br136_falseOut_ready;
  wire [6:0] buffer60_outs;
  wire  buffer60_outs_valid;
  wire  buffer60_outs_ready;
  wire [6:0] buffer61_outs;
  wire  buffer61_outs_valid;
  wire  buffer61_outs_ready;
  wire [6:0] cond_br137_trueOut;
  wire  cond_br137_trueOut_valid;
  wire  cond_br137_trueOut_ready;
  wire [6:0] cond_br137_falseOut;
  wire  cond_br137_falseOut_valid;
  wire  cond_br137_falseOut_ready;
  wire  cond_br138_trueOut_valid;
  wire  cond_br138_trueOut_ready;
  wire  cond_br138_falseOut_valid;
  wire  cond_br138_falseOut_ready;
  wire [4:0] cond_br139_trueOut;
  wire  cond_br139_trueOut_valid;
  wire  cond_br139_trueOut_ready;
  wire [4:0] cond_br139_falseOut;
  wire  cond_br139_falseOut_valid;
  wire  cond_br139_falseOut_ready;
  wire [4:0] buffer68_outs;
  wire  buffer68_outs_valid;
  wire  buffer68_outs_ready;
  wire [4:0] buffer69_outs;
  wire  buffer69_outs_valid;
  wire  buffer69_outs_ready;
  wire [4:0] fork37_outs_0;
  wire  fork37_outs_0_valid;
  wire  fork37_outs_0_ready;
  wire [4:0] fork37_outs_1;
  wire  fork37_outs_1_valid;
  wire  fork37_outs_1_ready;
  wire  buffer70_outs_valid;
  wire  buffer70_outs_ready;
  wire  buffer71_outs_valid;
  wire  buffer71_outs_ready;
  wire  fork38_outs_0_valid;
  wire  fork38_outs_0_ready;
  wire  fork38_outs_1_valid;
  wire  fork38_outs_1_ready;
  wire  fork38_outs_2_valid;
  wire  fork38_outs_2_ready;
  wire  fork38_outs_3_valid;
  wire  fork38_outs_3_ready;
  wire  fork38_outs_4_valid;
  wire  fork38_outs_4_ready;
  wire  fork38_outs_5_valid;
  wire  fork38_outs_5_ready;
  wire  fork38_outs_6_valid;
  wire  fork38_outs_6_ready;
  wire [36:0] constant307_outs;
  wire  constant307_outs_valid;
  wire  constant307_outs_ready;
  wire [30:0] constant497_outs;
  wire  constant497_outs_valid;
  wire  constant497_outs_ready;
  wire [26:0] constant309_outs;
  wire  constant309_outs_valid;
  wire  constant309_outs_ready;
  wire [20:0] constant498_outs;
  wire  constant498_outs_valid;
  wire  constant498_outs_ready;
  wire [16:0] constant311_outs;
  wire  constant311_outs_valid;
  wire  constant311_outs_ready;
  wire [11:0] constant312_outs;
  wire  constant312_outs_valid;
  wire  constant312_outs_ready;
  wire  source13_outs_valid;
  wire  source13_outs_ready;
  wire [4:0] constant499_outs;
  wire  constant499_outs_valid;
  wire  constant499_outs_ready;
  wire [0:0] cmpi12_result;
  wire  cmpi12_result_valid;
  wire  cmpi12_result_ready;
  wire [0:0] fork39_outs_0;
  wire  fork39_outs_0_valid;
  wire  fork39_outs_0_ready;
  wire [0:0] fork39_outs_1;
  wire  fork39_outs_1_valid;
  wire  fork39_outs_1_ready;
  wire [0:0] fork39_outs_2;
  wire  fork39_outs_2_valid;
  wire  fork39_outs_2_ready;
  wire [0:0] fork39_outs_3;
  wire  fork39_outs_3_valid;
  wire  fork39_outs_3_ready;
  wire [0:0] fork39_outs_4;
  wire  fork39_outs_4_valid;
  wire  fork39_outs_4_ready;
  wire [0:0] fork39_outs_5;
  wire  fork39_outs_5_valid;
  wire  fork39_outs_5_ready;
  wire [0:0] fork39_outs_6;
  wire  fork39_outs_6_valid;
  wire  fork39_outs_6_ready;
  wire [0:0] fork39_outs_7;
  wire  fork39_outs_7_valid;
  wire  fork39_outs_7_ready;
  wire [0:0] fork39_outs_8;
  wire  fork39_outs_8_valid;
  wire  fork39_outs_8_ready;
  wire [36:0] cond_br140_trueOut;
  wire  cond_br140_trueOut_valid;
  wire  cond_br140_trueOut_ready;
  wire [36:0] cond_br140_falseOut;
  wire  cond_br140_falseOut_valid;
  wire  cond_br140_falseOut_ready;
  wire [30:0] cond_br141_trueOut;
  wire  cond_br141_trueOut_valid;
  wire  cond_br141_trueOut_ready;
  wire [30:0] cond_br141_falseOut;
  wire  cond_br141_falseOut_valid;
  wire  cond_br141_falseOut_ready;
  wire [32:0] extsi174_outs;
  wire  extsi174_outs_valid;
  wire  extsi174_outs_ready;
  wire [26:0] cond_br142_trueOut;
  wire  cond_br142_trueOut_valid;
  wire  cond_br142_trueOut_ready;
  wire [26:0] cond_br142_falseOut;
  wire  cond_br142_falseOut_valid;
  wire  cond_br142_falseOut_ready;
  wire [20:0] cond_br143_trueOut;
  wire  cond_br143_trueOut_valid;
  wire  cond_br143_trueOut_ready;
  wire [20:0] cond_br143_falseOut;
  wire  cond_br143_falseOut_valid;
  wire  cond_br143_falseOut_ready;
  wire [21:0] extsi175_outs;
  wire  extsi175_outs_valid;
  wire  extsi175_outs_ready;
  wire [16:0] cond_br144_trueOut;
  wire  cond_br144_trueOut_valid;
  wire  cond_br144_trueOut_ready;
  wire [16:0] cond_br144_falseOut;
  wire  cond_br144_falseOut_valid;
  wire  cond_br144_falseOut_ready;
  wire [11:0] cond_br145_trueOut;
  wire  cond_br145_trueOut_valid;
  wire  cond_br145_trueOut_ready;
  wire [11:0] cond_br145_falseOut;
  wire  cond_br145_falseOut_valid;
  wire  cond_br145_falseOut_ready;
  wire [6:0] buffer66_outs;
  wire  buffer66_outs_valid;
  wire  buffer66_outs_ready;
  wire [6:0] buffer67_outs;
  wire  buffer67_outs_valid;
  wire  buffer67_outs_ready;
  wire [6:0] cond_br146_trueOut;
  wire  cond_br146_trueOut_valid;
  wire  cond_br146_trueOut_ready;
  wire [6:0] cond_br146_falseOut;
  wire  cond_br146_falseOut_valid;
  wire  cond_br146_falseOut_ready;
  wire  cond_br147_trueOut_valid;
  wire  cond_br147_trueOut_ready;
  wire  cond_br147_falseOut_valid;
  wire  cond_br147_falseOut_ready;
  wire [4:0] cond_br148_trueOut;
  wire  cond_br148_trueOut_valid;
  wire  cond_br148_trueOut_ready;
  wire [4:0] cond_br148_falseOut;
  wire  cond_br148_falseOut_valid;
  wire  cond_br148_falseOut_ready;
  wire [4:0] buffer74_outs;
  wire  buffer74_outs_valid;
  wire  buffer74_outs_ready;
  wire [4:0] buffer75_outs;
  wire  buffer75_outs_valid;
  wire  buffer75_outs_ready;
  wire [4:0] fork40_outs_0;
  wire  fork40_outs_0_valid;
  wire  fork40_outs_0_ready;
  wire [4:0] fork40_outs_1;
  wire  fork40_outs_1_valid;
  wire  fork40_outs_1_ready;
  wire  buffer76_outs_valid;
  wire  buffer76_outs_ready;
  wire  buffer77_outs_valid;
  wire  buffer77_outs_ready;
  wire  fork41_outs_0_valid;
  wire  fork41_outs_0_ready;
  wire  fork41_outs_1_valid;
  wire  fork41_outs_1_ready;
  wire  fork41_outs_2_valid;
  wire  fork41_outs_2_ready;
  wire  fork41_outs_3_valid;
  wire  fork41_outs_3_ready;
  wire  fork41_outs_4_valid;
  wire  fork41_outs_4_ready;
  wire  fork41_outs_5_valid;
  wire  fork41_outs_5_ready;
  wire  fork41_outs_6_valid;
  wire  fork41_outs_6_ready;
  wire [36:0] constant314_outs;
  wire  constant314_outs_valid;
  wire  constant314_outs_ready;
  wire [30:0] constant500_outs;
  wire  constant500_outs_valid;
  wire  constant500_outs_ready;
  wire [26:0] constant316_outs;
  wire  constant316_outs_valid;
  wire  constant316_outs_ready;
  wire [20:0] constant501_outs;
  wire  constant501_outs_valid;
  wire  constant501_outs_ready;
  wire [16:0] constant318_outs;
  wire  constant318_outs_valid;
  wire  constant318_outs_ready;
  wire [11:0] constant319_outs;
  wire  constant319_outs_valid;
  wire  constant319_outs_ready;
  wire  source14_outs_valid;
  wire  source14_outs_ready;
  wire [4:0] constant502_outs;
  wire  constant502_outs_valid;
  wire  constant502_outs_ready;
  wire [0:0] cmpi13_result;
  wire  cmpi13_result_valid;
  wire  cmpi13_result_ready;
  wire [0:0] fork42_outs_0;
  wire  fork42_outs_0_valid;
  wire  fork42_outs_0_ready;
  wire [0:0] fork42_outs_1;
  wire  fork42_outs_1_valid;
  wire  fork42_outs_1_ready;
  wire [0:0] fork42_outs_2;
  wire  fork42_outs_2_valid;
  wire  fork42_outs_2_ready;
  wire [0:0] fork42_outs_3;
  wire  fork42_outs_3_valid;
  wire  fork42_outs_3_ready;
  wire [0:0] fork42_outs_4;
  wire  fork42_outs_4_valid;
  wire  fork42_outs_4_ready;
  wire [0:0] fork42_outs_5;
  wire  fork42_outs_5_valid;
  wire  fork42_outs_5_ready;
  wire [0:0] fork42_outs_6;
  wire  fork42_outs_6_valid;
  wire  fork42_outs_6_ready;
  wire [0:0] fork42_outs_7;
  wire  fork42_outs_7_valid;
  wire  fork42_outs_7_ready;
  wire [0:0] fork42_outs_8;
  wire  fork42_outs_8_valid;
  wire  fork42_outs_8_ready;
  wire [36:0] cond_br149_trueOut;
  wire  cond_br149_trueOut_valid;
  wire  cond_br149_trueOut_ready;
  wire [36:0] cond_br149_falseOut;
  wire  cond_br149_falseOut_valid;
  wire  cond_br149_falseOut_ready;
  wire [30:0] cond_br150_trueOut;
  wire  cond_br150_trueOut_valid;
  wire  cond_br150_trueOut_ready;
  wire [30:0] cond_br150_falseOut;
  wire  cond_br150_falseOut_valid;
  wire  cond_br150_falseOut_ready;
  wire [32:0] extsi176_outs;
  wire  extsi176_outs_valid;
  wire  extsi176_outs_ready;
  wire [26:0] cond_br151_trueOut;
  wire  cond_br151_trueOut_valid;
  wire  cond_br151_trueOut_ready;
  wire [26:0] cond_br151_falseOut;
  wire  cond_br151_falseOut_valid;
  wire  cond_br151_falseOut_ready;
  wire [20:0] cond_br152_trueOut;
  wire  cond_br152_trueOut_valid;
  wire  cond_br152_trueOut_ready;
  wire [20:0] cond_br152_falseOut;
  wire  cond_br152_falseOut_valid;
  wire  cond_br152_falseOut_ready;
  wire [21:0] extsi177_outs;
  wire  extsi177_outs_valid;
  wire  extsi177_outs_ready;
  wire [16:0] cond_br153_trueOut;
  wire  cond_br153_trueOut_valid;
  wire  cond_br153_trueOut_ready;
  wire [16:0] cond_br153_falseOut;
  wire  cond_br153_falseOut_valid;
  wire  cond_br153_falseOut_ready;
  wire [11:0] cond_br154_trueOut;
  wire  cond_br154_trueOut_valid;
  wire  cond_br154_trueOut_ready;
  wire [11:0] cond_br154_falseOut;
  wire  cond_br154_falseOut_valid;
  wire  cond_br154_falseOut_ready;
  wire [6:0] buffer72_outs;
  wire  buffer72_outs_valid;
  wire  buffer72_outs_ready;
  wire [6:0] buffer73_outs;
  wire  buffer73_outs_valid;
  wire  buffer73_outs_ready;
  wire [6:0] cond_br155_trueOut;
  wire  cond_br155_trueOut_valid;
  wire  cond_br155_trueOut_ready;
  wire [6:0] cond_br155_falseOut;
  wire  cond_br155_falseOut_valid;
  wire  cond_br155_falseOut_ready;
  wire  cond_br156_trueOut_valid;
  wire  cond_br156_trueOut_ready;
  wire  cond_br156_falseOut_valid;
  wire  cond_br156_falseOut_ready;
  wire [4:0] cond_br157_trueOut;
  wire  cond_br157_trueOut_valid;
  wire  cond_br157_trueOut_ready;
  wire [4:0] cond_br157_falseOut;
  wire  cond_br157_falseOut_valid;
  wire  cond_br157_falseOut_ready;
  wire [4:0] buffer80_outs;
  wire  buffer80_outs_valid;
  wire  buffer80_outs_ready;
  wire [4:0] buffer81_outs;
  wire  buffer81_outs_valid;
  wire  buffer81_outs_ready;
  wire [4:0] fork43_outs_0;
  wire  fork43_outs_0_valid;
  wire  fork43_outs_0_ready;
  wire [4:0] fork43_outs_1;
  wire  fork43_outs_1_valid;
  wire  fork43_outs_1_ready;
  wire  buffer82_outs_valid;
  wire  buffer82_outs_ready;
  wire  buffer83_outs_valid;
  wire  buffer83_outs_ready;
  wire  fork44_outs_0_valid;
  wire  fork44_outs_0_ready;
  wire  fork44_outs_1_valid;
  wire  fork44_outs_1_ready;
  wire  fork44_outs_2_valid;
  wire  fork44_outs_2_ready;
  wire  fork44_outs_3_valid;
  wire  fork44_outs_3_ready;
  wire  fork44_outs_4_valid;
  wire  fork44_outs_4_ready;
  wire  fork44_outs_5_valid;
  wire  fork44_outs_5_ready;
  wire  fork44_outs_6_valid;
  wire  fork44_outs_6_ready;
  wire [36:0] constant321_outs;
  wire  constant321_outs_valid;
  wire  constant321_outs_ready;
  wire [30:0] constant503_outs;
  wire  constant503_outs_valid;
  wire  constant503_outs_ready;
  wire [26:0] constant323_outs;
  wire  constant323_outs_valid;
  wire  constant323_outs_ready;
  wire [20:0] constant504_outs;
  wire  constant504_outs_valid;
  wire  constant504_outs_ready;
  wire [16:0] constant325_outs;
  wire  constant325_outs_valid;
  wire  constant325_outs_ready;
  wire [11:0] constant326_outs;
  wire  constant326_outs_valid;
  wire  constant326_outs_ready;
  wire  source15_outs_valid;
  wire  source15_outs_ready;
  wire [4:0] constant505_outs;
  wire  constant505_outs_valid;
  wire  constant505_outs_ready;
  wire [0:0] cmpi14_result;
  wire  cmpi14_result_valid;
  wire  cmpi14_result_ready;
  wire [0:0] fork45_outs_0;
  wire  fork45_outs_0_valid;
  wire  fork45_outs_0_ready;
  wire [0:0] fork45_outs_1;
  wire  fork45_outs_1_valid;
  wire  fork45_outs_1_ready;
  wire [0:0] fork45_outs_2;
  wire  fork45_outs_2_valid;
  wire  fork45_outs_2_ready;
  wire [0:0] fork45_outs_3;
  wire  fork45_outs_3_valid;
  wire  fork45_outs_3_ready;
  wire [0:0] fork45_outs_4;
  wire  fork45_outs_4_valid;
  wire  fork45_outs_4_ready;
  wire [0:0] fork45_outs_5;
  wire  fork45_outs_5_valid;
  wire  fork45_outs_5_ready;
  wire [0:0] fork45_outs_6;
  wire  fork45_outs_6_valid;
  wire  fork45_outs_6_ready;
  wire [0:0] fork45_outs_7;
  wire  fork45_outs_7_valid;
  wire  fork45_outs_7_ready;
  wire [0:0] fork45_outs_8;
  wire  fork45_outs_8_valid;
  wire  fork45_outs_8_ready;
  wire [36:0] cond_br158_trueOut;
  wire  cond_br158_trueOut_valid;
  wire  cond_br158_trueOut_ready;
  wire [36:0] cond_br158_falseOut;
  wire  cond_br158_falseOut_valid;
  wire  cond_br158_falseOut_ready;
  wire [30:0] cond_br159_trueOut;
  wire  cond_br159_trueOut_valid;
  wire  cond_br159_trueOut_ready;
  wire [30:0] cond_br159_falseOut;
  wire  cond_br159_falseOut_valid;
  wire  cond_br159_falseOut_ready;
  wire [32:0] extsi178_outs;
  wire  extsi178_outs_valid;
  wire  extsi178_outs_ready;
  wire [26:0] cond_br160_trueOut;
  wire  cond_br160_trueOut_valid;
  wire  cond_br160_trueOut_ready;
  wire [26:0] cond_br160_falseOut;
  wire  cond_br160_falseOut_valid;
  wire  cond_br160_falseOut_ready;
  wire [20:0] cond_br161_trueOut;
  wire  cond_br161_trueOut_valid;
  wire  cond_br161_trueOut_ready;
  wire [20:0] cond_br161_falseOut;
  wire  cond_br161_falseOut_valid;
  wire  cond_br161_falseOut_ready;
  wire [21:0] extsi179_outs;
  wire  extsi179_outs_valid;
  wire  extsi179_outs_ready;
  wire [16:0] cond_br162_trueOut;
  wire  cond_br162_trueOut_valid;
  wire  cond_br162_trueOut_ready;
  wire [16:0] cond_br162_falseOut;
  wire  cond_br162_falseOut_valid;
  wire  cond_br162_falseOut_ready;
  wire [11:0] cond_br163_trueOut;
  wire  cond_br163_trueOut_valid;
  wire  cond_br163_trueOut_ready;
  wire [11:0] cond_br163_falseOut;
  wire  cond_br163_falseOut_valid;
  wire  cond_br163_falseOut_ready;
  wire [6:0] buffer78_outs;
  wire  buffer78_outs_valid;
  wire  buffer78_outs_ready;
  wire [6:0] buffer79_outs;
  wire  buffer79_outs_valid;
  wire  buffer79_outs_ready;
  wire [6:0] cond_br164_trueOut;
  wire  cond_br164_trueOut_valid;
  wire  cond_br164_trueOut_ready;
  wire [6:0] cond_br164_falseOut;
  wire  cond_br164_falseOut_valid;
  wire  cond_br164_falseOut_ready;
  wire  cond_br165_trueOut_valid;
  wire  cond_br165_trueOut_ready;
  wire  cond_br165_falseOut_valid;
  wire  cond_br165_falseOut_ready;
  wire [4:0] cond_br166_trueOut;
  wire  cond_br166_trueOut_valid;
  wire  cond_br166_trueOut_ready;
  wire [4:0] cond_br166_falseOut;
  wire  cond_br166_falseOut_valid;
  wire  cond_br166_falseOut_ready;
  wire [4:0] buffer86_outs;
  wire  buffer86_outs_valid;
  wire  buffer86_outs_ready;
  wire [4:0] buffer87_outs;
  wire  buffer87_outs_valid;
  wire  buffer87_outs_ready;
  wire [4:0] fork46_outs_0;
  wire  fork46_outs_0_valid;
  wire  fork46_outs_0_ready;
  wire [4:0] fork46_outs_1;
  wire  fork46_outs_1_valid;
  wire  fork46_outs_1_ready;
  wire  buffer88_outs_valid;
  wire  buffer88_outs_ready;
  wire  buffer89_outs_valid;
  wire  buffer89_outs_ready;
  wire  fork47_outs_0_valid;
  wire  fork47_outs_0_ready;
  wire  fork47_outs_1_valid;
  wire  fork47_outs_1_ready;
  wire  fork47_outs_2_valid;
  wire  fork47_outs_2_ready;
  wire  fork47_outs_3_valid;
  wire  fork47_outs_3_ready;
  wire  fork47_outs_4_valid;
  wire  fork47_outs_4_ready;
  wire  fork47_outs_5_valid;
  wire  fork47_outs_5_ready;
  wire  fork47_outs_6_valid;
  wire  fork47_outs_6_ready;
  wire [36:0] constant328_outs;
  wire  constant328_outs_valid;
  wire  constant328_outs_ready;
  wire [30:0] constant506_outs;
  wire  constant506_outs_valid;
  wire  constant506_outs_ready;
  wire [26:0] constant330_outs;
  wire  constant330_outs_valid;
  wire  constant330_outs_ready;
  wire [20:0] constant507_outs;
  wire  constant507_outs_valid;
  wire  constant507_outs_ready;
  wire [16:0] constant332_outs;
  wire  constant332_outs_valid;
  wire  constant332_outs_ready;
  wire [11:0] constant333_outs;
  wire  constant333_outs_valid;
  wire  constant333_outs_ready;
  wire  source16_outs_valid;
  wire  source16_outs_ready;
  wire [4:0] constant508_outs;
  wire  constant508_outs_valid;
  wire  constant508_outs_ready;
  wire [0:0] cmpi15_result;
  wire  cmpi15_result_valid;
  wire  cmpi15_result_ready;
  wire [0:0] fork48_outs_0;
  wire  fork48_outs_0_valid;
  wire  fork48_outs_0_ready;
  wire [0:0] fork48_outs_1;
  wire  fork48_outs_1_valid;
  wire  fork48_outs_1_ready;
  wire [0:0] fork48_outs_2;
  wire  fork48_outs_2_valid;
  wire  fork48_outs_2_ready;
  wire [0:0] fork48_outs_3;
  wire  fork48_outs_3_valid;
  wire  fork48_outs_3_ready;
  wire [0:0] fork48_outs_4;
  wire  fork48_outs_4_valid;
  wire  fork48_outs_4_ready;
  wire [0:0] fork48_outs_5;
  wire  fork48_outs_5_valid;
  wire  fork48_outs_5_ready;
  wire [0:0] fork48_outs_6;
  wire  fork48_outs_6_valid;
  wire  fork48_outs_6_ready;
  wire [0:0] fork48_outs_7;
  wire  fork48_outs_7_valid;
  wire  fork48_outs_7_ready;
  wire [0:0] fork48_outs_8;
  wire  fork48_outs_8_valid;
  wire  fork48_outs_8_ready;
  wire [36:0] cond_br167_trueOut;
  wire  cond_br167_trueOut_valid;
  wire  cond_br167_trueOut_ready;
  wire [36:0] cond_br167_falseOut;
  wire  cond_br167_falseOut_valid;
  wire  cond_br167_falseOut_ready;
  wire [30:0] cond_br168_trueOut;
  wire  cond_br168_trueOut_valid;
  wire  cond_br168_trueOut_ready;
  wire [30:0] cond_br168_falseOut;
  wire  cond_br168_falseOut_valid;
  wire  cond_br168_falseOut_ready;
  wire [32:0] extsi180_outs;
  wire  extsi180_outs_valid;
  wire  extsi180_outs_ready;
  wire [26:0] cond_br169_trueOut;
  wire  cond_br169_trueOut_valid;
  wire  cond_br169_trueOut_ready;
  wire [26:0] cond_br169_falseOut;
  wire  cond_br169_falseOut_valid;
  wire  cond_br169_falseOut_ready;
  wire [20:0] cond_br170_trueOut;
  wire  cond_br170_trueOut_valid;
  wire  cond_br170_trueOut_ready;
  wire [20:0] cond_br170_falseOut;
  wire  cond_br170_falseOut_valid;
  wire  cond_br170_falseOut_ready;
  wire [21:0] extsi181_outs;
  wire  extsi181_outs_valid;
  wire  extsi181_outs_ready;
  wire [16:0] cond_br171_trueOut;
  wire  cond_br171_trueOut_valid;
  wire  cond_br171_trueOut_ready;
  wire [16:0] cond_br171_falseOut;
  wire  cond_br171_falseOut_valid;
  wire  cond_br171_falseOut_ready;
  wire [11:0] cond_br172_trueOut;
  wire  cond_br172_trueOut_valid;
  wire  cond_br172_trueOut_ready;
  wire [11:0] cond_br172_falseOut;
  wire  cond_br172_falseOut_valid;
  wire  cond_br172_falseOut_ready;
  wire [6:0] buffer84_outs;
  wire  buffer84_outs_valid;
  wire  buffer84_outs_ready;
  wire [6:0] buffer85_outs;
  wire  buffer85_outs_valid;
  wire  buffer85_outs_ready;
  wire [6:0] cond_br173_trueOut;
  wire  cond_br173_trueOut_valid;
  wire  cond_br173_trueOut_ready;
  wire [6:0] cond_br173_falseOut;
  wire  cond_br173_falseOut_valid;
  wire  cond_br173_falseOut_ready;
  wire  cond_br174_trueOut_valid;
  wire  cond_br174_trueOut_ready;
  wire  cond_br174_falseOut_valid;
  wire  cond_br174_falseOut_ready;
  wire [4:0] cond_br175_trueOut;
  wire  cond_br175_trueOut_valid;
  wire  cond_br175_trueOut_ready;
  wire [4:0] cond_br175_falseOut;
  wire  cond_br175_falseOut_valid;
  wire  cond_br175_falseOut_ready;
  wire [4:0] buffer92_outs;
  wire  buffer92_outs_valid;
  wire  buffer92_outs_ready;
  wire [4:0] buffer93_outs;
  wire  buffer93_outs_valid;
  wire  buffer93_outs_ready;
  wire [4:0] fork49_outs_0;
  wire  fork49_outs_0_valid;
  wire  fork49_outs_0_ready;
  wire [4:0] fork49_outs_1;
  wire  fork49_outs_1_valid;
  wire  fork49_outs_1_ready;
  wire [5:0] extsi182_outs;
  wire  extsi182_outs_valid;
  wire  extsi182_outs_ready;
  wire  buffer94_outs_valid;
  wire  buffer94_outs_ready;
  wire  buffer95_outs_valid;
  wire  buffer95_outs_ready;
  wire  fork50_outs_0_valid;
  wire  fork50_outs_0_ready;
  wire  fork50_outs_1_valid;
  wire  fork50_outs_1_ready;
  wire  fork50_outs_2_valid;
  wire  fork50_outs_2_ready;
  wire  fork50_outs_3_valid;
  wire  fork50_outs_3_ready;
  wire  fork50_outs_4_valid;
  wire  fork50_outs_4_ready;
  wire  fork50_outs_5_valid;
  wire  fork50_outs_5_ready;
  wire  fork50_outs_6_valid;
  wire  fork50_outs_6_ready;
  wire [36:0] constant335_outs;
  wire  constant335_outs_valid;
  wire  constant335_outs_ready;
  wire [29:0] constant509_outs;
  wire  constant509_outs_valid;
  wire  constant509_outs_ready;
  wire [26:0] constant337_outs;
  wire  constant337_outs_valid;
  wire  constant337_outs_ready;
  wire [19:0] constant510_outs;
  wire  constant510_outs_valid;
  wire  constant510_outs_ready;
  wire [16:0] constant339_outs;
  wire  constant339_outs_valid;
  wire  constant339_outs_ready;
  wire [11:0] constant340_outs;
  wire  constant340_outs_valid;
  wire  constant340_outs_ready;
  wire  source17_outs_valid;
  wire  source17_outs_ready;
  wire [5:0] constant511_outs;
  wire  constant511_outs_valid;
  wire  constant511_outs_ready;
  wire [0:0] cmpi16_result;
  wire  cmpi16_result_valid;
  wire  cmpi16_result_ready;
  wire [0:0] fork51_outs_0;
  wire  fork51_outs_0_valid;
  wire  fork51_outs_0_ready;
  wire [0:0] fork51_outs_1;
  wire  fork51_outs_1_valid;
  wire  fork51_outs_1_ready;
  wire [0:0] fork51_outs_2;
  wire  fork51_outs_2_valid;
  wire  fork51_outs_2_ready;
  wire [0:0] fork51_outs_3;
  wire  fork51_outs_3_valid;
  wire  fork51_outs_3_ready;
  wire [0:0] fork51_outs_4;
  wire  fork51_outs_4_valid;
  wire  fork51_outs_4_ready;
  wire [0:0] fork51_outs_5;
  wire  fork51_outs_5_valid;
  wire  fork51_outs_5_ready;
  wire [0:0] fork51_outs_6;
  wire  fork51_outs_6_valid;
  wire  fork51_outs_6_ready;
  wire [0:0] fork51_outs_7;
  wire  fork51_outs_7_valid;
  wire  fork51_outs_7_ready;
  wire [0:0] fork51_outs_8;
  wire  fork51_outs_8_valid;
  wire  fork51_outs_8_ready;
  wire [36:0] cond_br176_trueOut;
  wire  cond_br176_trueOut_valid;
  wire  cond_br176_trueOut_ready;
  wire [36:0] cond_br176_falseOut;
  wire  cond_br176_falseOut_valid;
  wire  cond_br176_falseOut_ready;
  wire [29:0] cond_br177_trueOut;
  wire  cond_br177_trueOut_valid;
  wire  cond_br177_trueOut_ready;
  wire [29:0] cond_br177_falseOut;
  wire  cond_br177_falseOut_valid;
  wire  cond_br177_falseOut_ready;
  wire [32:0] extsi183_outs;
  wire  extsi183_outs_valid;
  wire  extsi183_outs_ready;
  wire [26:0] cond_br178_trueOut;
  wire  cond_br178_trueOut_valid;
  wire  cond_br178_trueOut_ready;
  wire [26:0] cond_br178_falseOut;
  wire  cond_br178_falseOut_valid;
  wire  cond_br178_falseOut_ready;
  wire [19:0] cond_br179_trueOut;
  wire  cond_br179_trueOut_valid;
  wire  cond_br179_trueOut_ready;
  wire [19:0] cond_br179_falseOut;
  wire  cond_br179_falseOut_valid;
  wire  cond_br179_falseOut_ready;
  wire [21:0] extsi184_outs;
  wire  extsi184_outs_valid;
  wire  extsi184_outs_ready;
  wire [16:0] cond_br180_trueOut;
  wire  cond_br180_trueOut_valid;
  wire  cond_br180_trueOut_ready;
  wire [16:0] cond_br180_falseOut;
  wire  cond_br180_falseOut_valid;
  wire  cond_br180_falseOut_ready;
  wire [11:0] cond_br181_trueOut;
  wire  cond_br181_trueOut_valid;
  wire  cond_br181_trueOut_ready;
  wire [11:0] cond_br181_falseOut;
  wire  cond_br181_falseOut_valid;
  wire  cond_br181_falseOut_ready;
  wire [6:0] buffer90_outs;
  wire  buffer90_outs_valid;
  wire  buffer90_outs_ready;
  wire [6:0] buffer91_outs;
  wire  buffer91_outs_valid;
  wire  buffer91_outs_ready;
  wire [6:0] cond_br182_trueOut;
  wire  cond_br182_trueOut_valid;
  wire  cond_br182_trueOut_ready;
  wire [6:0] cond_br182_falseOut;
  wire  cond_br182_falseOut_valid;
  wire  cond_br182_falseOut_ready;
  wire  cond_br183_trueOut_valid;
  wire  cond_br183_trueOut_ready;
  wire  cond_br183_falseOut_valid;
  wire  cond_br183_falseOut_ready;
  wire [4:0] cond_br184_trueOut;
  wire  cond_br184_trueOut_valid;
  wire  cond_br184_trueOut_ready;
  wire [4:0] cond_br184_falseOut;
  wire  cond_br184_falseOut_valid;
  wire  cond_br184_falseOut_ready;
  wire [4:0] buffer98_outs;
  wire  buffer98_outs_valid;
  wire  buffer98_outs_ready;
  wire [4:0] buffer99_outs;
  wire  buffer99_outs_valid;
  wire  buffer99_outs_ready;
  wire [4:0] fork52_outs_0;
  wire  fork52_outs_0_valid;
  wire  fork52_outs_0_ready;
  wire [4:0] fork52_outs_1;
  wire  fork52_outs_1_valid;
  wire  fork52_outs_1_ready;
  wire [5:0] extsi185_outs;
  wire  extsi185_outs_valid;
  wire  extsi185_outs_ready;
  wire  buffer100_outs_valid;
  wire  buffer100_outs_ready;
  wire  buffer101_outs_valid;
  wire  buffer101_outs_ready;
  wire  fork53_outs_0_valid;
  wire  fork53_outs_0_ready;
  wire  fork53_outs_1_valid;
  wire  fork53_outs_1_ready;
  wire  fork53_outs_2_valid;
  wire  fork53_outs_2_ready;
  wire  fork53_outs_3_valid;
  wire  fork53_outs_3_ready;
  wire  fork53_outs_4_valid;
  wire  fork53_outs_4_ready;
  wire  fork53_outs_5_valid;
  wire  fork53_outs_5_ready;
  wire  fork53_outs_6_valid;
  wire  fork53_outs_6_ready;
  wire [36:0] constant342_outs;
  wire  constant342_outs_valid;
  wire  constant342_outs_ready;
  wire [29:0] constant512_outs;
  wire  constant512_outs_valid;
  wire  constant512_outs_ready;
  wire [26:0] constant344_outs;
  wire  constant344_outs_valid;
  wire  constant344_outs_ready;
  wire [19:0] constant513_outs;
  wire  constant513_outs_valid;
  wire  constant513_outs_ready;
  wire [16:0] constant346_outs;
  wire  constant346_outs_valid;
  wire  constant346_outs_ready;
  wire [5:0] constant514_outs;
  wire  constant514_outs_valid;
  wire  constant514_outs_ready;
  wire  source18_outs_valid;
  wire  source18_outs_ready;
  wire [5:0] constant515_outs;
  wire  constant515_outs_valid;
  wire  constant515_outs_ready;
  wire [0:0] cmpi17_result;
  wire  cmpi17_result_valid;
  wire  cmpi17_result_ready;
  wire [0:0] fork54_outs_0;
  wire  fork54_outs_0_valid;
  wire  fork54_outs_0_ready;
  wire [0:0] fork54_outs_1;
  wire  fork54_outs_1_valid;
  wire  fork54_outs_1_ready;
  wire [0:0] fork54_outs_2;
  wire  fork54_outs_2_valid;
  wire  fork54_outs_2_ready;
  wire [0:0] fork54_outs_3;
  wire  fork54_outs_3_valid;
  wire  fork54_outs_3_ready;
  wire [0:0] fork54_outs_4;
  wire  fork54_outs_4_valid;
  wire  fork54_outs_4_ready;
  wire [0:0] fork54_outs_5;
  wire  fork54_outs_5_valid;
  wire  fork54_outs_5_ready;
  wire [0:0] fork54_outs_6;
  wire  fork54_outs_6_valid;
  wire  fork54_outs_6_ready;
  wire [0:0] fork54_outs_7;
  wire  fork54_outs_7_valid;
  wire  fork54_outs_7_ready;
  wire [0:0] fork54_outs_8;
  wire  fork54_outs_8_valid;
  wire  fork54_outs_8_ready;
  wire [36:0] cond_br185_trueOut;
  wire  cond_br185_trueOut_valid;
  wire  cond_br185_trueOut_ready;
  wire [36:0] cond_br185_falseOut;
  wire  cond_br185_falseOut_valid;
  wire  cond_br185_falseOut_ready;
  wire [29:0] cond_br186_trueOut;
  wire  cond_br186_trueOut_valid;
  wire  cond_br186_trueOut_ready;
  wire [29:0] cond_br186_falseOut;
  wire  cond_br186_falseOut_valid;
  wire  cond_br186_falseOut_ready;
  wire [32:0] extsi186_outs;
  wire  extsi186_outs_valid;
  wire  extsi186_outs_ready;
  wire [26:0] cond_br187_trueOut;
  wire  cond_br187_trueOut_valid;
  wire  cond_br187_trueOut_ready;
  wire [26:0] cond_br187_falseOut;
  wire  cond_br187_falseOut_valid;
  wire  cond_br187_falseOut_ready;
  wire [19:0] cond_br188_trueOut;
  wire  cond_br188_trueOut_valid;
  wire  cond_br188_trueOut_ready;
  wire [19:0] cond_br188_falseOut;
  wire  cond_br188_falseOut_valid;
  wire  cond_br188_falseOut_ready;
  wire [21:0] extsi187_outs;
  wire  extsi187_outs_valid;
  wire  extsi187_outs_ready;
  wire [16:0] cond_br189_trueOut;
  wire  cond_br189_trueOut_valid;
  wire  cond_br189_trueOut_ready;
  wire [16:0] cond_br189_falseOut;
  wire  cond_br189_falseOut_valid;
  wire  cond_br189_falseOut_ready;
  wire [5:0] cond_br190_trueOut;
  wire  cond_br190_trueOut_valid;
  wire  cond_br190_trueOut_ready;
  wire [5:0] cond_br190_falseOut;
  wire  cond_br190_falseOut_valid;
  wire  cond_br190_falseOut_ready;
  wire [11:0] extsi188_outs;
  wire  extsi188_outs_valid;
  wire  extsi188_outs_ready;
  wire [6:0] buffer96_outs;
  wire  buffer96_outs_valid;
  wire  buffer96_outs_ready;
  wire [6:0] buffer97_outs;
  wire  buffer97_outs_valid;
  wire  buffer97_outs_ready;
  wire [6:0] cond_br191_trueOut;
  wire  cond_br191_trueOut_valid;
  wire  cond_br191_trueOut_ready;
  wire [6:0] cond_br191_falseOut;
  wire  cond_br191_falseOut_valid;
  wire  cond_br191_falseOut_ready;
  wire  cond_br192_trueOut_valid;
  wire  cond_br192_trueOut_ready;
  wire  cond_br192_falseOut_valid;
  wire  cond_br192_falseOut_ready;
  wire [4:0] cond_br193_trueOut;
  wire  cond_br193_trueOut_valid;
  wire  cond_br193_trueOut_ready;
  wire [4:0] cond_br193_falseOut;
  wire  cond_br193_falseOut_valid;
  wire  cond_br193_falseOut_ready;
  wire [4:0] buffer104_outs;
  wire  buffer104_outs_valid;
  wire  buffer104_outs_ready;
  wire [4:0] buffer105_outs;
  wire  buffer105_outs_valid;
  wire  buffer105_outs_ready;
  wire [4:0] fork55_outs_0;
  wire  fork55_outs_0_valid;
  wire  fork55_outs_0_ready;
  wire [4:0] fork55_outs_1;
  wire  fork55_outs_1_valid;
  wire  fork55_outs_1_ready;
  wire [5:0] extsi189_outs;
  wire  extsi189_outs_valid;
  wire  extsi189_outs_ready;
  wire  buffer106_outs_valid;
  wire  buffer106_outs_ready;
  wire  buffer107_outs_valid;
  wire  buffer107_outs_ready;
  wire  fork56_outs_0_valid;
  wire  fork56_outs_0_ready;
  wire  fork56_outs_1_valid;
  wire  fork56_outs_1_ready;
  wire  fork56_outs_2_valid;
  wire  fork56_outs_2_ready;
  wire  fork56_outs_3_valid;
  wire  fork56_outs_3_ready;
  wire  fork56_outs_4_valid;
  wire  fork56_outs_4_ready;
  wire  fork56_outs_5_valid;
  wire  fork56_outs_5_ready;
  wire  fork56_outs_6_valid;
  wire  fork56_outs_6_ready;
  wire [36:0] constant349_outs;
  wire  constant349_outs_valid;
  wire  constant349_outs_ready;
  wire [29:0] constant516_outs;
  wire  constant516_outs_valid;
  wire  constant516_outs_ready;
  wire [26:0] constant351_outs;
  wire  constant351_outs_valid;
  wire  constant351_outs_ready;
  wire [19:0] constant517_outs;
  wire  constant517_outs_valid;
  wire  constant517_outs_ready;
  wire [16:0] constant353_outs;
  wire  constant353_outs_valid;
  wire  constant353_outs_ready;
  wire [6:0] constant518_outs;
  wire  constant518_outs_valid;
  wire  constant518_outs_ready;
  wire  source19_outs_valid;
  wire  source19_outs_ready;
  wire [5:0] constant519_outs;
  wire  constant519_outs_valid;
  wire  constant519_outs_ready;
  wire [0:0] cmpi18_result;
  wire  cmpi18_result_valid;
  wire  cmpi18_result_ready;
  wire [0:0] fork57_outs_0;
  wire  fork57_outs_0_valid;
  wire  fork57_outs_0_ready;
  wire [0:0] fork57_outs_1;
  wire  fork57_outs_1_valid;
  wire  fork57_outs_1_ready;
  wire [0:0] fork57_outs_2;
  wire  fork57_outs_2_valid;
  wire  fork57_outs_2_ready;
  wire [0:0] fork57_outs_3;
  wire  fork57_outs_3_valid;
  wire  fork57_outs_3_ready;
  wire [0:0] fork57_outs_4;
  wire  fork57_outs_4_valid;
  wire  fork57_outs_4_ready;
  wire [0:0] fork57_outs_5;
  wire  fork57_outs_5_valid;
  wire  fork57_outs_5_ready;
  wire [0:0] fork57_outs_6;
  wire  fork57_outs_6_valid;
  wire  fork57_outs_6_ready;
  wire [0:0] fork57_outs_7;
  wire  fork57_outs_7_valid;
  wire  fork57_outs_7_ready;
  wire [0:0] fork57_outs_8;
  wire  fork57_outs_8_valid;
  wire  fork57_outs_8_ready;
  wire [36:0] cond_br194_trueOut;
  wire  cond_br194_trueOut_valid;
  wire  cond_br194_trueOut_ready;
  wire [36:0] cond_br194_falseOut;
  wire  cond_br194_falseOut_valid;
  wire  cond_br194_falseOut_ready;
  wire [29:0] cond_br195_trueOut;
  wire  cond_br195_trueOut_valid;
  wire  cond_br195_trueOut_ready;
  wire [29:0] cond_br195_falseOut;
  wire  cond_br195_falseOut_valid;
  wire  cond_br195_falseOut_ready;
  wire [32:0] extsi190_outs;
  wire  extsi190_outs_valid;
  wire  extsi190_outs_ready;
  wire [26:0] cond_br196_trueOut;
  wire  cond_br196_trueOut_valid;
  wire  cond_br196_trueOut_ready;
  wire [26:0] cond_br196_falseOut;
  wire  cond_br196_falseOut_valid;
  wire  cond_br196_falseOut_ready;
  wire [19:0] cond_br197_trueOut;
  wire  cond_br197_trueOut_valid;
  wire  cond_br197_trueOut_ready;
  wire [19:0] cond_br197_falseOut;
  wire  cond_br197_falseOut_valid;
  wire  cond_br197_falseOut_ready;
  wire [21:0] extsi191_outs;
  wire  extsi191_outs_valid;
  wire  extsi191_outs_ready;
  wire [16:0] cond_br198_trueOut;
  wire  cond_br198_trueOut_valid;
  wire  cond_br198_trueOut_ready;
  wire [16:0] cond_br198_falseOut;
  wire  cond_br198_falseOut_valid;
  wire  cond_br198_falseOut_ready;
  wire [6:0] cond_br199_trueOut;
  wire  cond_br199_trueOut_valid;
  wire  cond_br199_trueOut_ready;
  wire [6:0] cond_br199_falseOut;
  wire  cond_br199_falseOut_valid;
  wire  cond_br199_falseOut_ready;
  wire [11:0] extsi192_outs;
  wire  extsi192_outs_valid;
  wire  extsi192_outs_ready;
  wire [6:0] buffer102_outs;
  wire  buffer102_outs_valid;
  wire  buffer102_outs_ready;
  wire [6:0] buffer103_outs;
  wire  buffer103_outs_valid;
  wire  buffer103_outs_ready;
  wire [6:0] cond_br200_trueOut;
  wire  cond_br200_trueOut_valid;
  wire  cond_br200_trueOut_ready;
  wire [6:0] cond_br200_falseOut;
  wire  cond_br200_falseOut_valid;
  wire  cond_br200_falseOut_ready;
  wire  cond_br201_trueOut_valid;
  wire  cond_br201_trueOut_ready;
  wire  cond_br201_falseOut_valid;
  wire  cond_br201_falseOut_ready;
  wire [4:0] cond_br202_trueOut;
  wire  cond_br202_trueOut_valid;
  wire  cond_br202_trueOut_ready;
  wire [4:0] cond_br202_falseOut;
  wire  cond_br202_falseOut_valid;
  wire  cond_br202_falseOut_ready;
  wire [4:0] buffer110_outs;
  wire  buffer110_outs_valid;
  wire  buffer110_outs_ready;
  wire [4:0] buffer111_outs;
  wire  buffer111_outs_valid;
  wire  buffer111_outs_ready;
  wire [4:0] fork58_outs_0;
  wire  fork58_outs_0_valid;
  wire  fork58_outs_0_ready;
  wire [4:0] fork58_outs_1;
  wire  fork58_outs_1_valid;
  wire  fork58_outs_1_ready;
  wire [5:0] extsi193_outs;
  wire  extsi193_outs_valid;
  wire  extsi193_outs_ready;
  wire  buffer112_outs_valid;
  wire  buffer112_outs_ready;
  wire  buffer113_outs_valid;
  wire  buffer113_outs_ready;
  wire  fork59_outs_0_valid;
  wire  fork59_outs_0_ready;
  wire  fork59_outs_1_valid;
  wire  fork59_outs_1_ready;
  wire  fork59_outs_2_valid;
  wire  fork59_outs_2_ready;
  wire  fork59_outs_3_valid;
  wire  fork59_outs_3_ready;
  wire  fork59_outs_4_valid;
  wire  fork59_outs_4_ready;
  wire  fork59_outs_5_valid;
  wire  fork59_outs_5_ready;
  wire  fork59_outs_6_valid;
  wire  fork59_outs_6_ready;
  wire [36:0] constant356_outs;
  wire  constant356_outs_valid;
  wire  constant356_outs_ready;
  wire [29:0] constant520_outs;
  wire  constant520_outs_valid;
  wire  constant520_outs_ready;
  wire [26:0] constant358_outs;
  wire  constant358_outs_valid;
  wire  constant358_outs_ready;
  wire [19:0] constant521_outs;
  wire  constant521_outs_valid;
  wire  constant521_outs_ready;
  wire [16:0] constant360_outs;
  wire  constant360_outs_valid;
  wire  constant360_outs_ready;
  wire [6:0] constant522_outs;
  wire  constant522_outs_valid;
  wire  constant522_outs_ready;
  wire  source20_outs_valid;
  wire  source20_outs_ready;
  wire [5:0] constant523_outs;
  wire  constant523_outs_valid;
  wire  constant523_outs_ready;
  wire [0:0] cmpi19_result;
  wire  cmpi19_result_valid;
  wire  cmpi19_result_ready;
  wire [0:0] fork60_outs_0;
  wire  fork60_outs_0_valid;
  wire  fork60_outs_0_ready;
  wire [0:0] fork60_outs_1;
  wire  fork60_outs_1_valid;
  wire  fork60_outs_1_ready;
  wire [0:0] fork60_outs_2;
  wire  fork60_outs_2_valid;
  wire  fork60_outs_2_ready;
  wire [0:0] fork60_outs_3;
  wire  fork60_outs_3_valid;
  wire  fork60_outs_3_ready;
  wire [0:0] fork60_outs_4;
  wire  fork60_outs_4_valid;
  wire  fork60_outs_4_ready;
  wire [0:0] fork60_outs_5;
  wire  fork60_outs_5_valid;
  wire  fork60_outs_5_ready;
  wire [0:0] fork60_outs_6;
  wire  fork60_outs_6_valid;
  wire  fork60_outs_6_ready;
  wire [0:0] fork60_outs_7;
  wire  fork60_outs_7_valid;
  wire  fork60_outs_7_ready;
  wire [0:0] fork60_outs_8;
  wire  fork60_outs_8_valid;
  wire  fork60_outs_8_ready;
  wire [36:0] cond_br203_trueOut;
  wire  cond_br203_trueOut_valid;
  wire  cond_br203_trueOut_ready;
  wire [36:0] cond_br203_falseOut;
  wire  cond_br203_falseOut_valid;
  wire  cond_br203_falseOut_ready;
  wire [29:0] cond_br204_trueOut;
  wire  cond_br204_trueOut_valid;
  wire  cond_br204_trueOut_ready;
  wire [29:0] cond_br204_falseOut;
  wire  cond_br204_falseOut_valid;
  wire  cond_br204_falseOut_ready;
  wire [32:0] extsi194_outs;
  wire  extsi194_outs_valid;
  wire  extsi194_outs_ready;
  wire [26:0] cond_br205_trueOut;
  wire  cond_br205_trueOut_valid;
  wire  cond_br205_trueOut_ready;
  wire [26:0] cond_br205_falseOut;
  wire  cond_br205_falseOut_valid;
  wire  cond_br205_falseOut_ready;
  wire [19:0] cond_br206_trueOut;
  wire  cond_br206_trueOut_valid;
  wire  cond_br206_trueOut_ready;
  wire [19:0] cond_br206_falseOut;
  wire  cond_br206_falseOut_valid;
  wire  cond_br206_falseOut_ready;
  wire [21:0] extsi195_outs;
  wire  extsi195_outs_valid;
  wire  extsi195_outs_ready;
  wire [16:0] cond_br207_trueOut;
  wire  cond_br207_trueOut_valid;
  wire  cond_br207_trueOut_ready;
  wire [16:0] cond_br207_falseOut;
  wire  cond_br207_falseOut_valid;
  wire  cond_br207_falseOut_ready;
  wire [6:0] cond_br208_trueOut;
  wire  cond_br208_trueOut_valid;
  wire  cond_br208_trueOut_ready;
  wire [6:0] cond_br208_falseOut;
  wire  cond_br208_falseOut_valid;
  wire  cond_br208_falseOut_ready;
  wire [11:0] extsi196_outs;
  wire  extsi196_outs_valid;
  wire  extsi196_outs_ready;
  wire [6:0] buffer108_outs;
  wire  buffer108_outs_valid;
  wire  buffer108_outs_ready;
  wire [6:0] buffer109_outs;
  wire  buffer109_outs_valid;
  wire  buffer109_outs_ready;
  wire [6:0] cond_br209_trueOut;
  wire  cond_br209_trueOut_valid;
  wire  cond_br209_trueOut_ready;
  wire [6:0] cond_br209_falseOut;
  wire  cond_br209_falseOut_valid;
  wire  cond_br209_falseOut_ready;
  wire  cond_br210_trueOut_valid;
  wire  cond_br210_trueOut_ready;
  wire  cond_br210_falseOut_valid;
  wire  cond_br210_falseOut_ready;
  wire [4:0] cond_br211_trueOut;
  wire  cond_br211_trueOut_valid;
  wire  cond_br211_trueOut_ready;
  wire [4:0] cond_br211_falseOut;
  wire  cond_br211_falseOut_valid;
  wire  cond_br211_falseOut_ready;
  wire [4:0] buffer116_outs;
  wire  buffer116_outs_valid;
  wire  buffer116_outs_ready;
  wire [4:0] buffer117_outs;
  wire  buffer117_outs_valid;
  wire  buffer117_outs_ready;
  wire [4:0] fork61_outs_0;
  wire  fork61_outs_0_valid;
  wire  fork61_outs_0_ready;
  wire [4:0] fork61_outs_1;
  wire  fork61_outs_1_valid;
  wire  fork61_outs_1_ready;
  wire [5:0] extsi197_outs;
  wire  extsi197_outs_valid;
  wire  extsi197_outs_ready;
  wire  buffer118_outs_valid;
  wire  buffer118_outs_ready;
  wire  buffer119_outs_valid;
  wire  buffer119_outs_ready;
  wire  fork62_outs_0_valid;
  wire  fork62_outs_0_ready;
  wire  fork62_outs_1_valid;
  wire  fork62_outs_1_ready;
  wire  fork62_outs_2_valid;
  wire  fork62_outs_2_ready;
  wire  fork62_outs_3_valid;
  wire  fork62_outs_3_ready;
  wire  fork62_outs_4_valid;
  wire  fork62_outs_4_ready;
  wire  fork62_outs_5_valid;
  wire  fork62_outs_5_ready;
  wire  fork62_outs_6_valid;
  wire  fork62_outs_6_ready;
  wire [36:0] constant363_outs;
  wire  constant363_outs_valid;
  wire  constant363_outs_ready;
  wire [28:0] constant524_outs;
  wire  constant524_outs_valid;
  wire  constant524_outs_ready;
  wire [26:0] constant365_outs;
  wire  constant365_outs_valid;
  wire  constant365_outs_ready;
  wire [19:0] constant525_outs;
  wire  constant525_outs_valid;
  wire  constant525_outs_ready;
  wire [16:0] constant367_outs;
  wire  constant367_outs_valid;
  wire  constant367_outs_ready;
  wire [6:0] constant526_outs;
  wire  constant526_outs_valid;
  wire  constant526_outs_ready;
  wire  source21_outs_valid;
  wire  source21_outs_ready;
  wire [5:0] constant527_outs;
  wire  constant527_outs_valid;
  wire  constant527_outs_ready;
  wire [0:0] cmpi20_result;
  wire  cmpi20_result_valid;
  wire  cmpi20_result_ready;
  wire [0:0] fork63_outs_0;
  wire  fork63_outs_0_valid;
  wire  fork63_outs_0_ready;
  wire [0:0] fork63_outs_1;
  wire  fork63_outs_1_valid;
  wire  fork63_outs_1_ready;
  wire [0:0] fork63_outs_2;
  wire  fork63_outs_2_valid;
  wire  fork63_outs_2_ready;
  wire [0:0] fork63_outs_3;
  wire  fork63_outs_3_valid;
  wire  fork63_outs_3_ready;
  wire [0:0] fork63_outs_4;
  wire  fork63_outs_4_valid;
  wire  fork63_outs_4_ready;
  wire [0:0] fork63_outs_5;
  wire  fork63_outs_5_valid;
  wire  fork63_outs_5_ready;
  wire [0:0] fork63_outs_6;
  wire  fork63_outs_6_valid;
  wire  fork63_outs_6_ready;
  wire [0:0] fork63_outs_7;
  wire  fork63_outs_7_valid;
  wire  fork63_outs_7_ready;
  wire [0:0] fork63_outs_8;
  wire  fork63_outs_8_valid;
  wire  fork63_outs_8_ready;
  wire [36:0] cond_br212_trueOut;
  wire  cond_br212_trueOut_valid;
  wire  cond_br212_trueOut_ready;
  wire [36:0] cond_br212_falseOut;
  wire  cond_br212_falseOut_valid;
  wire  cond_br212_falseOut_ready;
  wire [28:0] cond_br213_trueOut;
  wire  cond_br213_trueOut_valid;
  wire  cond_br213_trueOut_ready;
  wire [28:0] cond_br213_falseOut;
  wire  cond_br213_falseOut_valid;
  wire  cond_br213_falseOut_ready;
  wire [32:0] extsi198_outs;
  wire  extsi198_outs_valid;
  wire  extsi198_outs_ready;
  wire [26:0] cond_br214_trueOut;
  wire  cond_br214_trueOut_valid;
  wire  cond_br214_trueOut_ready;
  wire [26:0] cond_br214_falseOut;
  wire  cond_br214_falseOut_valid;
  wire  cond_br214_falseOut_ready;
  wire [19:0] cond_br215_trueOut;
  wire  cond_br215_trueOut_valid;
  wire  cond_br215_trueOut_ready;
  wire [19:0] cond_br215_falseOut;
  wire  cond_br215_falseOut_valid;
  wire  cond_br215_falseOut_ready;
  wire [21:0] extsi199_outs;
  wire  extsi199_outs_valid;
  wire  extsi199_outs_ready;
  wire [16:0] cond_br216_trueOut;
  wire  cond_br216_trueOut_valid;
  wire  cond_br216_trueOut_ready;
  wire [16:0] cond_br216_falseOut;
  wire  cond_br216_falseOut_valid;
  wire  cond_br216_falseOut_ready;
  wire [6:0] cond_br217_trueOut;
  wire  cond_br217_trueOut_valid;
  wire  cond_br217_trueOut_ready;
  wire [6:0] cond_br217_falseOut;
  wire  cond_br217_falseOut_valid;
  wire  cond_br217_falseOut_ready;
  wire [11:0] extsi200_outs;
  wire  extsi200_outs_valid;
  wire  extsi200_outs_ready;
  wire [6:0] buffer114_outs;
  wire  buffer114_outs_valid;
  wire  buffer114_outs_ready;
  wire [6:0] buffer115_outs;
  wire  buffer115_outs_valid;
  wire  buffer115_outs_ready;
  wire [6:0] cond_br218_trueOut;
  wire  cond_br218_trueOut_valid;
  wire  cond_br218_trueOut_ready;
  wire [6:0] cond_br218_falseOut;
  wire  cond_br218_falseOut_valid;
  wire  cond_br218_falseOut_ready;
  wire  cond_br219_trueOut_valid;
  wire  cond_br219_trueOut_ready;
  wire  cond_br219_falseOut_valid;
  wire  cond_br219_falseOut_ready;
  wire [4:0] cond_br220_trueOut;
  wire  cond_br220_trueOut_valid;
  wire  cond_br220_trueOut_ready;
  wire [4:0] cond_br220_falseOut;
  wire  cond_br220_falseOut_valid;
  wire  cond_br220_falseOut_ready;
  wire [4:0] buffer122_outs;
  wire  buffer122_outs_valid;
  wire  buffer122_outs_ready;
  wire [4:0] buffer123_outs;
  wire  buffer123_outs_valid;
  wire  buffer123_outs_ready;
  wire [4:0] fork64_outs_0;
  wire  fork64_outs_0_valid;
  wire  fork64_outs_0_ready;
  wire [4:0] fork64_outs_1;
  wire  fork64_outs_1_valid;
  wire  fork64_outs_1_ready;
  wire [5:0] extsi201_outs;
  wire  extsi201_outs_valid;
  wire  extsi201_outs_ready;
  wire  buffer124_outs_valid;
  wire  buffer124_outs_ready;
  wire  buffer125_outs_valid;
  wire  buffer125_outs_ready;
  wire  fork65_outs_0_valid;
  wire  fork65_outs_0_ready;
  wire  fork65_outs_1_valid;
  wire  fork65_outs_1_ready;
  wire  fork65_outs_2_valid;
  wire  fork65_outs_2_ready;
  wire  fork65_outs_3_valid;
  wire  fork65_outs_3_ready;
  wire  fork65_outs_4_valid;
  wire  fork65_outs_4_ready;
  wire  fork65_outs_5_valid;
  wire  fork65_outs_5_ready;
  wire  fork65_outs_6_valid;
  wire  fork65_outs_6_ready;
  wire [36:0] constant370_outs;
  wire  constant370_outs_valid;
  wire  constant370_outs_ready;
  wire [28:0] constant528_outs;
  wire  constant528_outs_valid;
  wire  constant528_outs_ready;
  wire [26:0] constant372_outs;
  wire  constant372_outs_valid;
  wire  constant372_outs_ready;
  wire [18:0] constant529_outs;
  wire  constant529_outs_valid;
  wire  constant529_outs_ready;
  wire [16:0] constant374_outs;
  wire  constant374_outs_valid;
  wire  constant374_outs_ready;
  wire [7:0] constant530_outs;
  wire  constant530_outs_valid;
  wire  constant530_outs_ready;
  wire  source22_outs_valid;
  wire  source22_outs_ready;
  wire [5:0] constant531_outs;
  wire  constant531_outs_valid;
  wire  constant531_outs_ready;
  wire [0:0] cmpi21_result;
  wire  cmpi21_result_valid;
  wire  cmpi21_result_ready;
  wire [0:0] fork66_outs_0;
  wire  fork66_outs_0_valid;
  wire  fork66_outs_0_ready;
  wire [0:0] fork66_outs_1;
  wire  fork66_outs_1_valid;
  wire  fork66_outs_1_ready;
  wire [0:0] fork66_outs_2;
  wire  fork66_outs_2_valid;
  wire  fork66_outs_2_ready;
  wire [0:0] fork66_outs_3;
  wire  fork66_outs_3_valid;
  wire  fork66_outs_3_ready;
  wire [0:0] fork66_outs_4;
  wire  fork66_outs_4_valid;
  wire  fork66_outs_4_ready;
  wire [0:0] fork66_outs_5;
  wire  fork66_outs_5_valid;
  wire  fork66_outs_5_ready;
  wire [0:0] fork66_outs_6;
  wire  fork66_outs_6_valid;
  wire  fork66_outs_6_ready;
  wire [0:0] fork66_outs_7;
  wire  fork66_outs_7_valid;
  wire  fork66_outs_7_ready;
  wire [0:0] fork66_outs_8;
  wire  fork66_outs_8_valid;
  wire  fork66_outs_8_ready;
  wire [36:0] cond_br221_trueOut;
  wire  cond_br221_trueOut_valid;
  wire  cond_br221_trueOut_ready;
  wire [36:0] cond_br221_falseOut;
  wire  cond_br221_falseOut_valid;
  wire  cond_br221_falseOut_ready;
  wire [28:0] cond_br222_trueOut;
  wire  cond_br222_trueOut_valid;
  wire  cond_br222_trueOut_ready;
  wire [28:0] cond_br222_falseOut;
  wire  cond_br222_falseOut_valid;
  wire  cond_br222_falseOut_ready;
  wire [32:0] extsi202_outs;
  wire  extsi202_outs_valid;
  wire  extsi202_outs_ready;
  wire [26:0] cond_br223_trueOut;
  wire  cond_br223_trueOut_valid;
  wire  cond_br223_trueOut_ready;
  wire [26:0] cond_br223_falseOut;
  wire  cond_br223_falseOut_valid;
  wire  cond_br223_falseOut_ready;
  wire [18:0] cond_br224_trueOut;
  wire  cond_br224_trueOut_valid;
  wire  cond_br224_trueOut_ready;
  wire [18:0] cond_br224_falseOut;
  wire  cond_br224_falseOut_valid;
  wire  cond_br224_falseOut_ready;
  wire [21:0] extsi203_outs;
  wire  extsi203_outs_valid;
  wire  extsi203_outs_ready;
  wire [16:0] cond_br225_trueOut;
  wire  cond_br225_trueOut_valid;
  wire  cond_br225_trueOut_ready;
  wire [16:0] cond_br225_falseOut;
  wire  cond_br225_falseOut_valid;
  wire  cond_br225_falseOut_ready;
  wire [7:0] cond_br226_trueOut;
  wire  cond_br226_trueOut_valid;
  wire  cond_br226_trueOut_ready;
  wire [7:0] cond_br226_falseOut;
  wire  cond_br226_falseOut_valid;
  wire  cond_br226_falseOut_ready;
  wire [11:0] extsi204_outs;
  wire  extsi204_outs_valid;
  wire  extsi204_outs_ready;
  wire [6:0] buffer120_outs;
  wire  buffer120_outs_valid;
  wire  buffer120_outs_ready;
  wire [6:0] buffer121_outs;
  wire  buffer121_outs_valid;
  wire  buffer121_outs_ready;
  wire [6:0] cond_br227_trueOut;
  wire  cond_br227_trueOut_valid;
  wire  cond_br227_trueOut_ready;
  wire [6:0] cond_br227_falseOut;
  wire  cond_br227_falseOut_valid;
  wire  cond_br227_falseOut_ready;
  wire  cond_br228_trueOut_valid;
  wire  cond_br228_trueOut_ready;
  wire  cond_br228_falseOut_valid;
  wire  cond_br228_falseOut_ready;
  wire [4:0] cond_br229_trueOut;
  wire  cond_br229_trueOut_valid;
  wire  cond_br229_trueOut_ready;
  wire [4:0] cond_br229_falseOut;
  wire  cond_br229_falseOut_valid;
  wire  cond_br229_falseOut_ready;
  wire [4:0] buffer128_outs;
  wire  buffer128_outs_valid;
  wire  buffer128_outs_ready;
  wire [4:0] buffer129_outs;
  wire  buffer129_outs_valid;
  wire  buffer129_outs_ready;
  wire [4:0] fork67_outs_0;
  wire  fork67_outs_0_valid;
  wire  fork67_outs_0_ready;
  wire [4:0] fork67_outs_1;
  wire  fork67_outs_1_valid;
  wire  fork67_outs_1_ready;
  wire [5:0] extsi205_outs;
  wire  extsi205_outs_valid;
  wire  extsi205_outs_ready;
  wire  buffer130_outs_valid;
  wire  buffer130_outs_ready;
  wire  buffer131_outs_valid;
  wire  buffer131_outs_ready;
  wire  fork68_outs_0_valid;
  wire  fork68_outs_0_ready;
  wire  fork68_outs_1_valid;
  wire  fork68_outs_1_ready;
  wire  fork68_outs_2_valid;
  wire  fork68_outs_2_ready;
  wire  fork68_outs_3_valid;
  wire  fork68_outs_3_ready;
  wire  fork68_outs_4_valid;
  wire  fork68_outs_4_ready;
  wire  fork68_outs_5_valid;
  wire  fork68_outs_5_ready;
  wire  fork68_outs_6_valid;
  wire  fork68_outs_6_ready;
  wire [36:0] constant377_outs;
  wire  constant377_outs_valid;
  wire  constant377_outs_ready;
  wire [28:0] constant532_outs;
  wire  constant532_outs_valid;
  wire  constant532_outs_ready;
  wire [26:0] constant379_outs;
  wire  constant379_outs_valid;
  wire  constant379_outs_ready;
  wire [18:0] constant533_outs;
  wire  constant533_outs_valid;
  wire  constant533_outs_ready;
  wire [16:0] constant381_outs;
  wire  constant381_outs_valid;
  wire  constant381_outs_ready;
  wire [6:0] constant534_outs;
  wire  constant534_outs_valid;
  wire  constant534_outs_ready;
  wire  source23_outs_valid;
  wire  source23_outs_ready;
  wire [5:0] constant535_outs;
  wire  constant535_outs_valid;
  wire  constant535_outs_ready;
  wire [0:0] cmpi22_result;
  wire  cmpi22_result_valid;
  wire  cmpi22_result_ready;
  wire [0:0] fork69_outs_0;
  wire  fork69_outs_0_valid;
  wire  fork69_outs_0_ready;
  wire [0:0] fork69_outs_1;
  wire  fork69_outs_1_valid;
  wire  fork69_outs_1_ready;
  wire [0:0] fork69_outs_2;
  wire  fork69_outs_2_valid;
  wire  fork69_outs_2_ready;
  wire [0:0] fork69_outs_3;
  wire  fork69_outs_3_valid;
  wire  fork69_outs_3_ready;
  wire [0:0] fork69_outs_4;
  wire  fork69_outs_4_valid;
  wire  fork69_outs_4_ready;
  wire [0:0] fork69_outs_5;
  wire  fork69_outs_5_valid;
  wire  fork69_outs_5_ready;
  wire [0:0] fork69_outs_6;
  wire  fork69_outs_6_valid;
  wire  fork69_outs_6_ready;
  wire [0:0] fork69_outs_7;
  wire  fork69_outs_7_valid;
  wire  fork69_outs_7_ready;
  wire [0:0] fork69_outs_8;
  wire  fork69_outs_8_valid;
  wire  fork69_outs_8_ready;
  wire [36:0] cond_br230_trueOut;
  wire  cond_br230_trueOut_valid;
  wire  cond_br230_trueOut_ready;
  wire [36:0] cond_br230_falseOut;
  wire  cond_br230_falseOut_valid;
  wire  cond_br230_falseOut_ready;
  wire [28:0] cond_br231_trueOut;
  wire  cond_br231_trueOut_valid;
  wire  cond_br231_trueOut_ready;
  wire [28:0] cond_br231_falseOut;
  wire  cond_br231_falseOut_valid;
  wire  cond_br231_falseOut_ready;
  wire [32:0] extsi206_outs;
  wire  extsi206_outs_valid;
  wire  extsi206_outs_ready;
  wire [26:0] cond_br232_trueOut;
  wire  cond_br232_trueOut_valid;
  wire  cond_br232_trueOut_ready;
  wire [26:0] cond_br232_falseOut;
  wire  cond_br232_falseOut_valid;
  wire  cond_br232_falseOut_ready;
  wire [18:0] cond_br233_trueOut;
  wire  cond_br233_trueOut_valid;
  wire  cond_br233_trueOut_ready;
  wire [18:0] cond_br233_falseOut;
  wire  cond_br233_falseOut_valid;
  wire  cond_br233_falseOut_ready;
  wire [21:0] extsi207_outs;
  wire  extsi207_outs_valid;
  wire  extsi207_outs_ready;
  wire [16:0] cond_br234_trueOut;
  wire  cond_br234_trueOut_valid;
  wire  cond_br234_trueOut_ready;
  wire [16:0] cond_br234_falseOut;
  wire  cond_br234_falseOut_valid;
  wire  cond_br234_falseOut_ready;
  wire [6:0] cond_br235_trueOut;
  wire  cond_br235_trueOut_valid;
  wire  cond_br235_trueOut_ready;
  wire [6:0] cond_br235_falseOut;
  wire  cond_br235_falseOut_valid;
  wire  cond_br235_falseOut_ready;
  wire [11:0] extsi208_outs;
  wire  extsi208_outs_valid;
  wire  extsi208_outs_ready;
  wire [6:0] buffer126_outs;
  wire  buffer126_outs_valid;
  wire  buffer126_outs_ready;
  wire [6:0] buffer127_outs;
  wire  buffer127_outs_valid;
  wire  buffer127_outs_ready;
  wire [6:0] cond_br236_trueOut;
  wire  cond_br236_trueOut_valid;
  wire  cond_br236_trueOut_ready;
  wire [6:0] cond_br236_falseOut;
  wire  cond_br236_falseOut_valid;
  wire  cond_br236_falseOut_ready;
  wire  cond_br237_trueOut_valid;
  wire  cond_br237_trueOut_ready;
  wire  cond_br237_falseOut_valid;
  wire  cond_br237_falseOut_ready;
  wire [4:0] cond_br238_trueOut;
  wire  cond_br238_trueOut_valid;
  wire  cond_br238_trueOut_ready;
  wire [4:0] cond_br238_falseOut;
  wire  cond_br238_falseOut_valid;
  wire  cond_br238_falseOut_ready;
  wire [4:0] buffer134_outs;
  wire  buffer134_outs_valid;
  wire  buffer134_outs_ready;
  wire [4:0] buffer135_outs;
  wire  buffer135_outs_valid;
  wire  buffer135_outs_ready;
  wire [4:0] fork70_outs_0;
  wire  fork70_outs_0_valid;
  wire  fork70_outs_0_ready;
  wire [4:0] fork70_outs_1;
  wire  fork70_outs_1_valid;
  wire  fork70_outs_1_ready;
  wire [5:0] extsi209_outs;
  wire  extsi209_outs_valid;
  wire  extsi209_outs_ready;
  wire  buffer136_outs_valid;
  wire  buffer136_outs_ready;
  wire  buffer137_outs_valid;
  wire  buffer137_outs_ready;
  wire  fork71_outs_0_valid;
  wire  fork71_outs_0_ready;
  wire  fork71_outs_1_valid;
  wire  fork71_outs_1_ready;
  wire  fork71_outs_2_valid;
  wire  fork71_outs_2_ready;
  wire  fork71_outs_3_valid;
  wire  fork71_outs_3_ready;
  wire  fork71_outs_4_valid;
  wire  fork71_outs_4_ready;
  wire  fork71_outs_5_valid;
  wire  fork71_outs_5_ready;
  wire  fork71_outs_6_valid;
  wire  fork71_outs_6_ready;
  wire [6:0] constant536_outs;
  wire  constant536_outs_valid;
  wire  constant536_outs_ready;
  wire [36:0] constant385_outs;
  wire  constant385_outs_valid;
  wire  constant385_outs_ready;
  wire [28:0] constant537_outs;
  wire  constant537_outs_valid;
  wire  constant537_outs_ready;
  wire [26:0] constant387_outs;
  wire  constant387_outs_valid;
  wire  constant387_outs_ready;
  wire [18:0] constant538_outs;
  wire  constant538_outs_valid;
  wire  constant538_outs_ready;
  wire [16:0] constant389_outs;
  wire  constant389_outs_valid;
  wire  constant389_outs_ready;
  wire  source24_outs_valid;
  wire  source24_outs_ready;
  wire [5:0] constant539_outs;
  wire  constant539_outs_valid;
  wire  constant539_outs_ready;
  wire [0:0] cmpi23_result;
  wire  cmpi23_result_valid;
  wire  cmpi23_result_ready;
  wire [0:0] fork72_outs_0;
  wire  fork72_outs_0_valid;
  wire  fork72_outs_0_ready;
  wire [0:0] fork72_outs_1;
  wire  fork72_outs_1_valid;
  wire  fork72_outs_1_ready;
  wire [0:0] fork72_outs_2;
  wire  fork72_outs_2_valid;
  wire  fork72_outs_2_ready;
  wire [0:0] fork72_outs_3;
  wire  fork72_outs_3_valid;
  wire  fork72_outs_3_ready;
  wire [0:0] fork72_outs_4;
  wire  fork72_outs_4_valid;
  wire  fork72_outs_4_ready;
  wire [0:0] fork72_outs_5;
  wire  fork72_outs_5_valid;
  wire  fork72_outs_5_ready;
  wire [0:0] fork72_outs_6;
  wire  fork72_outs_6_valid;
  wire  fork72_outs_6_ready;
  wire [0:0] fork72_outs_7;
  wire  fork72_outs_7_valid;
  wire  fork72_outs_7_ready;
  wire [0:0] fork72_outs_8;
  wire  fork72_outs_8_valid;
  wire  fork72_outs_8_ready;
  wire [36:0] cond_br239_trueOut;
  wire  cond_br239_trueOut_valid;
  wire  cond_br239_trueOut_ready;
  wire [36:0] cond_br239_falseOut;
  wire  cond_br239_falseOut_valid;
  wire  cond_br239_falseOut_ready;
  wire [28:0] cond_br240_trueOut;
  wire  cond_br240_trueOut_valid;
  wire  cond_br240_trueOut_ready;
  wire [28:0] cond_br240_falseOut;
  wire  cond_br240_falseOut_valid;
  wire  cond_br240_falseOut_ready;
  wire [32:0] extsi210_outs;
  wire  extsi210_outs_valid;
  wire  extsi210_outs_ready;
  wire [26:0] cond_br241_trueOut;
  wire  cond_br241_trueOut_valid;
  wire  cond_br241_trueOut_ready;
  wire [26:0] cond_br241_falseOut;
  wire  cond_br241_falseOut_valid;
  wire  cond_br241_falseOut_ready;
  wire [18:0] cond_br242_trueOut;
  wire  cond_br242_trueOut_valid;
  wire  cond_br242_trueOut_ready;
  wire [18:0] cond_br242_falseOut;
  wire  cond_br242_falseOut_valid;
  wire  cond_br242_falseOut_ready;
  wire [21:0] extsi211_outs;
  wire  extsi211_outs_valid;
  wire  extsi211_outs_ready;
  wire [16:0] cond_br243_trueOut;
  wire  cond_br243_trueOut_valid;
  wire  cond_br243_trueOut_ready;
  wire [16:0] cond_br243_falseOut;
  wire  cond_br243_falseOut_valid;
  wire  cond_br243_falseOut_ready;
  wire [6:0] cond_br244_trueOut;
  wire  cond_br244_trueOut_valid;
  wire  cond_br244_trueOut_ready;
  wire [6:0] cond_br244_falseOut;
  wire  cond_br244_falseOut_valid;
  wire  cond_br244_falseOut_ready;
  wire [11:0] extsi212_outs;
  wire  extsi212_outs_valid;
  wire  extsi212_outs_ready;
  wire [6:0] buffer132_outs;
  wire  buffer132_outs_valid;
  wire  buffer132_outs_ready;
  wire [6:0] buffer133_outs;
  wire  buffer133_outs_valid;
  wire  buffer133_outs_ready;
  wire [6:0] cond_br245_trueOut;
  wire  cond_br245_trueOut_valid;
  wire  cond_br245_trueOut_ready;
  wire [6:0] cond_br245_falseOut;
  wire  cond_br245_falseOut_valid;
  wire  cond_br245_falseOut_ready;
  wire  cond_br246_trueOut_valid;
  wire  cond_br246_trueOut_ready;
  wire  cond_br246_falseOut_valid;
  wire  cond_br246_falseOut_ready;
  wire [4:0] cond_br247_trueOut;
  wire  cond_br247_trueOut_valid;
  wire  cond_br247_trueOut_ready;
  wire [4:0] cond_br247_falseOut;
  wire  cond_br247_falseOut_valid;
  wire  cond_br247_falseOut_ready;
  wire [4:0] buffer140_outs;
  wire  buffer140_outs_valid;
  wire  buffer140_outs_ready;
  wire [4:0] buffer141_outs;
  wire  buffer141_outs_valid;
  wire  buffer141_outs_ready;
  wire [4:0] fork73_outs_0;
  wire  fork73_outs_0_valid;
  wire  fork73_outs_0_ready;
  wire [4:0] fork73_outs_1;
  wire  fork73_outs_1_valid;
  wire  fork73_outs_1_ready;
  wire [5:0] extsi213_outs;
  wire  extsi213_outs_valid;
  wire  extsi213_outs_ready;
  wire  buffer142_outs_valid;
  wire  buffer142_outs_ready;
  wire  buffer143_outs_valid;
  wire  buffer143_outs_ready;
  wire  fork74_outs_0_valid;
  wire  fork74_outs_0_ready;
  wire  fork74_outs_1_valid;
  wire  fork74_outs_1_ready;
  wire  fork74_outs_2_valid;
  wire  fork74_outs_2_ready;
  wire  fork74_outs_3_valid;
  wire  fork74_outs_3_ready;
  wire  fork74_outs_4_valid;
  wire  fork74_outs_4_ready;
  wire  fork74_outs_5_valid;
  wire  fork74_outs_5_ready;
  wire  fork74_outs_6_valid;
  wire  fork74_outs_6_ready;
  wire [36:0] constant391_outs;
  wire  constant391_outs_valid;
  wire  constant391_outs_ready;
  wire [27:0] constant540_outs;
  wire  constant540_outs_valid;
  wire  constant540_outs_ready;
  wire [26:0] constant393_outs;
  wire  constant393_outs_valid;
  wire  constant393_outs_ready;
  wire [18:0] constant541_outs;
  wire  constant541_outs_valid;
  wire  constant541_outs_ready;
  wire [16:0] constant395_outs;
  wire  constant395_outs_valid;
  wire  constant395_outs_ready;
  wire [6:0] constant542_outs;
  wire  constant542_outs_valid;
  wire  constant542_outs_ready;
  wire  source25_outs_valid;
  wire  source25_outs_ready;
  wire [5:0] constant543_outs;
  wire  constant543_outs_valid;
  wire  constant543_outs_ready;
  wire [0:0] cmpi24_result;
  wire  cmpi24_result_valid;
  wire  cmpi24_result_ready;
  wire [0:0] fork75_outs_0;
  wire  fork75_outs_0_valid;
  wire  fork75_outs_0_ready;
  wire [0:0] fork75_outs_1;
  wire  fork75_outs_1_valid;
  wire  fork75_outs_1_ready;
  wire [0:0] fork75_outs_2;
  wire  fork75_outs_2_valid;
  wire  fork75_outs_2_ready;
  wire [0:0] fork75_outs_3;
  wire  fork75_outs_3_valid;
  wire  fork75_outs_3_ready;
  wire [0:0] fork75_outs_4;
  wire  fork75_outs_4_valid;
  wire  fork75_outs_4_ready;
  wire [0:0] fork75_outs_5;
  wire  fork75_outs_5_valid;
  wire  fork75_outs_5_ready;
  wire [0:0] fork75_outs_6;
  wire  fork75_outs_6_valid;
  wire  fork75_outs_6_ready;
  wire [0:0] fork75_outs_7;
  wire  fork75_outs_7_valid;
  wire  fork75_outs_7_ready;
  wire [0:0] fork75_outs_8;
  wire  fork75_outs_8_valid;
  wire  fork75_outs_8_ready;
  wire [36:0] cond_br248_trueOut;
  wire  cond_br248_trueOut_valid;
  wire  cond_br248_trueOut_ready;
  wire [36:0] cond_br248_falseOut;
  wire  cond_br248_falseOut_valid;
  wire  cond_br248_falseOut_ready;
  wire [27:0] cond_br249_trueOut;
  wire  cond_br249_trueOut_valid;
  wire  cond_br249_trueOut_ready;
  wire [27:0] cond_br249_falseOut;
  wire  cond_br249_falseOut_valid;
  wire  cond_br249_falseOut_ready;
  wire [32:0] extsi214_outs;
  wire  extsi214_outs_valid;
  wire  extsi214_outs_ready;
  wire [26:0] cond_br250_trueOut;
  wire  cond_br250_trueOut_valid;
  wire  cond_br250_trueOut_ready;
  wire [26:0] cond_br250_falseOut;
  wire  cond_br250_falseOut_valid;
  wire  cond_br250_falseOut_ready;
  wire [18:0] cond_br251_trueOut;
  wire  cond_br251_trueOut_valid;
  wire  cond_br251_trueOut_ready;
  wire [18:0] cond_br251_falseOut;
  wire  cond_br251_falseOut_valid;
  wire  cond_br251_falseOut_ready;
  wire [21:0] extsi215_outs;
  wire  extsi215_outs_valid;
  wire  extsi215_outs_ready;
  wire [16:0] cond_br252_trueOut;
  wire  cond_br252_trueOut_valid;
  wire  cond_br252_trueOut_ready;
  wire [16:0] cond_br252_falseOut;
  wire  cond_br252_falseOut_valid;
  wire  cond_br252_falseOut_ready;
  wire [6:0] cond_br253_trueOut;
  wire  cond_br253_trueOut_valid;
  wire  cond_br253_trueOut_ready;
  wire [6:0] cond_br253_falseOut;
  wire  cond_br253_falseOut_valid;
  wire  cond_br253_falseOut_ready;
  wire [11:0] extsi216_outs;
  wire  extsi216_outs_valid;
  wire  extsi216_outs_ready;
  wire [6:0] buffer138_outs;
  wire  buffer138_outs_valid;
  wire  buffer138_outs_ready;
  wire [6:0] buffer139_outs;
  wire  buffer139_outs_valid;
  wire  buffer139_outs_ready;
  wire [6:0] cond_br254_trueOut;
  wire  cond_br254_trueOut_valid;
  wire  cond_br254_trueOut_ready;
  wire [6:0] cond_br254_falseOut;
  wire  cond_br254_falseOut_valid;
  wire  cond_br254_falseOut_ready;
  wire  cond_br255_trueOut_valid;
  wire  cond_br255_trueOut_ready;
  wire  cond_br255_falseOut_valid;
  wire  cond_br255_falseOut_ready;
  wire [4:0] cond_br256_trueOut;
  wire  cond_br256_trueOut_valid;
  wire  cond_br256_trueOut_ready;
  wire [4:0] cond_br256_falseOut;
  wire  cond_br256_falseOut_valid;
  wire  cond_br256_falseOut_ready;
  wire [4:0] buffer146_outs;
  wire  buffer146_outs_valid;
  wire  buffer146_outs_ready;
  wire [4:0] buffer147_outs;
  wire  buffer147_outs_valid;
  wire  buffer147_outs_ready;
  wire [4:0] fork76_outs_0;
  wire  fork76_outs_0_valid;
  wire  fork76_outs_0_ready;
  wire [4:0] fork76_outs_1;
  wire  fork76_outs_1_valid;
  wire  fork76_outs_1_ready;
  wire [5:0] extsi217_outs;
  wire  extsi217_outs_valid;
  wire  extsi217_outs_ready;
  wire  buffer148_outs_valid;
  wire  buffer148_outs_ready;
  wire  buffer149_outs_valid;
  wire  buffer149_outs_ready;
  wire  fork77_outs_0_valid;
  wire  fork77_outs_0_ready;
  wire  fork77_outs_1_valid;
  wire  fork77_outs_1_ready;
  wire  fork77_outs_2_valid;
  wire  fork77_outs_2_ready;
  wire  fork77_outs_3_valid;
  wire  fork77_outs_3_ready;
  wire  fork77_outs_4_valid;
  wire  fork77_outs_4_ready;
  wire  fork77_outs_5_valid;
  wire  fork77_outs_5_ready;
  wire  fork77_outs_6_valid;
  wire  fork77_outs_6_ready;
  wire [36:0] constant398_outs;
  wire  constant398_outs_valid;
  wire  constant398_outs_ready;
  wire [27:0] constant544_outs;
  wire  constant544_outs_valid;
  wire  constant544_outs_ready;
  wire [26:0] constant400_outs;
  wire  constant400_outs_valid;
  wire  constant400_outs_ready;
  wire [17:0] constant545_outs;
  wire  constant545_outs_valid;
  wire  constant545_outs_ready;
  wire [16:0] constant402_outs;
  wire  constant402_outs_valid;
  wire  constant402_outs_ready;
  wire [6:0] constant546_outs;
  wire  constant546_outs_valid;
  wire  constant546_outs_ready;
  wire  source26_outs_valid;
  wire  source26_outs_ready;
  wire [5:0] constant547_outs;
  wire  constant547_outs_valid;
  wire  constant547_outs_ready;
  wire [0:0] cmpi25_result;
  wire  cmpi25_result_valid;
  wire  cmpi25_result_ready;
  wire [0:0] fork78_outs_0;
  wire  fork78_outs_0_valid;
  wire  fork78_outs_0_ready;
  wire [0:0] fork78_outs_1;
  wire  fork78_outs_1_valid;
  wire  fork78_outs_1_ready;
  wire [0:0] fork78_outs_2;
  wire  fork78_outs_2_valid;
  wire  fork78_outs_2_ready;
  wire [0:0] fork78_outs_3;
  wire  fork78_outs_3_valid;
  wire  fork78_outs_3_ready;
  wire [0:0] fork78_outs_4;
  wire  fork78_outs_4_valid;
  wire  fork78_outs_4_ready;
  wire [0:0] fork78_outs_5;
  wire  fork78_outs_5_valid;
  wire  fork78_outs_5_ready;
  wire [0:0] fork78_outs_6;
  wire  fork78_outs_6_valid;
  wire  fork78_outs_6_ready;
  wire [0:0] fork78_outs_7;
  wire  fork78_outs_7_valid;
  wire  fork78_outs_7_ready;
  wire [0:0] fork78_outs_8;
  wire  fork78_outs_8_valid;
  wire  fork78_outs_8_ready;
  wire [36:0] cond_br257_trueOut;
  wire  cond_br257_trueOut_valid;
  wire  cond_br257_trueOut_ready;
  wire [36:0] cond_br257_falseOut;
  wire  cond_br257_falseOut_valid;
  wire  cond_br257_falseOut_ready;
  wire [27:0] cond_br258_trueOut;
  wire  cond_br258_trueOut_valid;
  wire  cond_br258_trueOut_ready;
  wire [27:0] cond_br258_falseOut;
  wire  cond_br258_falseOut_valid;
  wire  cond_br258_falseOut_ready;
  wire [32:0] extsi218_outs;
  wire  extsi218_outs_valid;
  wire  extsi218_outs_ready;
  wire [26:0] cond_br259_trueOut;
  wire  cond_br259_trueOut_valid;
  wire  cond_br259_trueOut_ready;
  wire [26:0] cond_br259_falseOut;
  wire  cond_br259_falseOut_valid;
  wire  cond_br259_falseOut_ready;
  wire [17:0] cond_br260_trueOut;
  wire  cond_br260_trueOut_valid;
  wire  cond_br260_trueOut_ready;
  wire [17:0] cond_br260_falseOut;
  wire  cond_br260_falseOut_valid;
  wire  cond_br260_falseOut_ready;
  wire [21:0] extsi219_outs;
  wire  extsi219_outs_valid;
  wire  extsi219_outs_ready;
  wire [16:0] cond_br261_trueOut;
  wire  cond_br261_trueOut_valid;
  wire  cond_br261_trueOut_ready;
  wire [16:0] cond_br261_falseOut;
  wire  cond_br261_falseOut_valid;
  wire  cond_br261_falseOut_ready;
  wire [6:0] cond_br262_trueOut;
  wire  cond_br262_trueOut_valid;
  wire  cond_br262_trueOut_ready;
  wire [6:0] cond_br262_falseOut;
  wire  cond_br262_falseOut_valid;
  wire  cond_br262_falseOut_ready;
  wire [11:0] extsi220_outs;
  wire  extsi220_outs_valid;
  wire  extsi220_outs_ready;
  wire [6:0] buffer144_outs;
  wire  buffer144_outs_valid;
  wire  buffer144_outs_ready;
  wire [6:0] buffer145_outs;
  wire  buffer145_outs_valid;
  wire  buffer145_outs_ready;
  wire [6:0] cond_br263_trueOut;
  wire  cond_br263_trueOut_valid;
  wire  cond_br263_trueOut_ready;
  wire [6:0] cond_br263_falseOut;
  wire  cond_br263_falseOut_valid;
  wire  cond_br263_falseOut_ready;
  wire  cond_br264_trueOut_valid;
  wire  cond_br264_trueOut_ready;
  wire  cond_br264_falseOut_valid;
  wire  cond_br264_falseOut_ready;
  wire [4:0] cond_br265_trueOut;
  wire  cond_br265_trueOut_valid;
  wire  cond_br265_trueOut_ready;
  wire [4:0] cond_br265_falseOut;
  wire  cond_br265_falseOut_valid;
  wire  cond_br265_falseOut_ready;
  wire [4:0] buffer152_outs;
  wire  buffer152_outs_valid;
  wire  buffer152_outs_ready;
  wire [4:0] buffer153_outs;
  wire  buffer153_outs_valid;
  wire  buffer153_outs_ready;
  wire [4:0] fork79_outs_0;
  wire  fork79_outs_0_valid;
  wire  fork79_outs_0_ready;
  wire [4:0] fork79_outs_1;
  wire  fork79_outs_1_valid;
  wire  fork79_outs_1_ready;
  wire [5:0] extsi221_outs;
  wire  extsi221_outs_valid;
  wire  extsi221_outs_ready;
  wire  buffer154_outs_valid;
  wire  buffer154_outs_ready;
  wire  buffer155_outs_valid;
  wire  buffer155_outs_ready;
  wire  fork80_outs_0_valid;
  wire  fork80_outs_0_ready;
  wire  fork80_outs_1_valid;
  wire  fork80_outs_1_ready;
  wire  fork80_outs_2_valid;
  wire  fork80_outs_2_ready;
  wire  fork80_outs_3_valid;
  wire  fork80_outs_3_ready;
  wire  fork80_outs_4_valid;
  wire  fork80_outs_4_ready;
  wire  fork80_outs_5_valid;
  wire  fork80_outs_5_ready;
  wire  fork80_outs_6_valid;
  wire  fork80_outs_6_ready;
  wire [36:0] constant405_outs;
  wire  constant405_outs_valid;
  wire  constant405_outs_ready;
  wire [27:0] constant548_outs;
  wire  constant548_outs_valid;
  wire  constant548_outs_ready;
  wire [26:0] constant407_outs;
  wire  constant407_outs_valid;
  wire  constant407_outs_ready;
  wire [17:0] constant549_outs;
  wire  constant549_outs_valid;
  wire  constant549_outs_ready;
  wire [16:0] constant409_outs;
  wire  constant409_outs_valid;
  wire  constant409_outs_ready;
  wire [6:0] constant550_outs;
  wire  constant550_outs_valid;
  wire  constant550_outs_ready;
  wire  source27_outs_valid;
  wire  source27_outs_ready;
  wire [5:0] constant551_outs;
  wire  constant551_outs_valid;
  wire  constant551_outs_ready;
  wire [0:0] cmpi26_result;
  wire  cmpi26_result_valid;
  wire  cmpi26_result_ready;
  wire [0:0] fork81_outs_0;
  wire  fork81_outs_0_valid;
  wire  fork81_outs_0_ready;
  wire [0:0] fork81_outs_1;
  wire  fork81_outs_1_valid;
  wire  fork81_outs_1_ready;
  wire [0:0] fork81_outs_2;
  wire  fork81_outs_2_valid;
  wire  fork81_outs_2_ready;
  wire [0:0] fork81_outs_3;
  wire  fork81_outs_3_valid;
  wire  fork81_outs_3_ready;
  wire [0:0] fork81_outs_4;
  wire  fork81_outs_4_valid;
  wire  fork81_outs_4_ready;
  wire [0:0] fork81_outs_5;
  wire  fork81_outs_5_valid;
  wire  fork81_outs_5_ready;
  wire [0:0] fork81_outs_6;
  wire  fork81_outs_6_valid;
  wire  fork81_outs_6_ready;
  wire [0:0] fork81_outs_7;
  wire  fork81_outs_7_valid;
  wire  fork81_outs_7_ready;
  wire [0:0] fork81_outs_8;
  wire  fork81_outs_8_valid;
  wire  fork81_outs_8_ready;
  wire [36:0] cond_br266_trueOut;
  wire  cond_br266_trueOut_valid;
  wire  cond_br266_trueOut_ready;
  wire [36:0] cond_br266_falseOut;
  wire  cond_br266_falseOut_valid;
  wire  cond_br266_falseOut_ready;
  wire [27:0] cond_br267_trueOut;
  wire  cond_br267_trueOut_valid;
  wire  cond_br267_trueOut_ready;
  wire [27:0] cond_br267_falseOut;
  wire  cond_br267_falseOut_valid;
  wire  cond_br267_falseOut_ready;
  wire [32:0] extsi222_outs;
  wire  extsi222_outs_valid;
  wire  extsi222_outs_ready;
  wire [26:0] cond_br268_trueOut;
  wire  cond_br268_trueOut_valid;
  wire  cond_br268_trueOut_ready;
  wire [26:0] cond_br268_falseOut;
  wire  cond_br268_falseOut_valid;
  wire  cond_br268_falseOut_ready;
  wire [17:0] cond_br269_trueOut;
  wire  cond_br269_trueOut_valid;
  wire  cond_br269_trueOut_ready;
  wire [17:0] cond_br269_falseOut;
  wire  cond_br269_falseOut_valid;
  wire  cond_br269_falseOut_ready;
  wire [21:0] extsi223_outs;
  wire  extsi223_outs_valid;
  wire  extsi223_outs_ready;
  wire [16:0] cond_br270_trueOut;
  wire  cond_br270_trueOut_valid;
  wire  cond_br270_trueOut_ready;
  wire [16:0] cond_br270_falseOut;
  wire  cond_br270_falseOut_valid;
  wire  cond_br270_falseOut_ready;
  wire [6:0] cond_br271_trueOut;
  wire  cond_br271_trueOut_valid;
  wire  cond_br271_trueOut_ready;
  wire [6:0] cond_br271_falseOut;
  wire  cond_br271_falseOut_valid;
  wire  cond_br271_falseOut_ready;
  wire [11:0] extsi224_outs;
  wire  extsi224_outs_valid;
  wire  extsi224_outs_ready;
  wire [6:0] buffer150_outs;
  wire  buffer150_outs_valid;
  wire  buffer150_outs_ready;
  wire [6:0] buffer151_outs;
  wire  buffer151_outs_valid;
  wire  buffer151_outs_ready;
  wire [6:0] cond_br272_trueOut;
  wire  cond_br272_trueOut_valid;
  wire  cond_br272_trueOut_ready;
  wire [6:0] cond_br272_falseOut;
  wire  cond_br272_falseOut_valid;
  wire  cond_br272_falseOut_ready;
  wire  cond_br273_trueOut_valid;
  wire  cond_br273_trueOut_ready;
  wire  cond_br273_falseOut_valid;
  wire  cond_br273_falseOut_ready;
  wire [4:0] cond_br274_trueOut;
  wire  cond_br274_trueOut_valid;
  wire  cond_br274_trueOut_ready;
  wire [4:0] cond_br274_falseOut;
  wire  cond_br274_falseOut_valid;
  wire  cond_br274_falseOut_ready;
  wire [4:0] buffer158_outs;
  wire  buffer158_outs_valid;
  wire  buffer158_outs_ready;
  wire [4:0] buffer159_outs;
  wire  buffer159_outs_valid;
  wire  buffer159_outs_ready;
  wire [4:0] fork82_outs_0;
  wire  fork82_outs_0_valid;
  wire  fork82_outs_0_ready;
  wire [4:0] fork82_outs_1;
  wire  fork82_outs_1_valid;
  wire  fork82_outs_1_ready;
  wire [5:0] extsi225_outs;
  wire  extsi225_outs_valid;
  wire  extsi225_outs_ready;
  wire  buffer160_outs_valid;
  wire  buffer160_outs_ready;
  wire  buffer161_outs_valid;
  wire  buffer161_outs_ready;
  wire  fork83_outs_0_valid;
  wire  fork83_outs_0_ready;
  wire  fork83_outs_1_valid;
  wire  fork83_outs_1_ready;
  wire  fork83_outs_2_valid;
  wire  fork83_outs_2_ready;
  wire  fork83_outs_3_valid;
  wire  fork83_outs_3_ready;
  wire  fork83_outs_4_valid;
  wire  fork83_outs_4_ready;
  wire  fork83_outs_5_valid;
  wire  fork83_outs_5_ready;
  wire  fork83_outs_6_valid;
  wire  fork83_outs_6_ready;
  wire [36:0] constant412_outs;
  wire  constant412_outs_valid;
  wire  constant412_outs_ready;
  wire [26:0] constant552_outs;
  wire  constant552_outs_valid;
  wire  constant552_outs_ready;
  wire [26:0] constant414_outs;
  wire  constant414_outs_valid;
  wire  constant414_outs_ready;
  wire [17:0] constant553_outs;
  wire  constant553_outs_valid;
  wire  constant553_outs_ready;
  wire [16:0] constant416_outs;
  wire  constant416_outs_valid;
  wire  constant416_outs_ready;
  wire [6:0] constant554_outs;
  wire  constant554_outs_valid;
  wire  constant554_outs_ready;
  wire  source28_outs_valid;
  wire  source28_outs_ready;
  wire [5:0] constant555_outs;
  wire  constant555_outs_valid;
  wire  constant555_outs_ready;
  wire [0:0] cmpi27_result;
  wire  cmpi27_result_valid;
  wire  cmpi27_result_ready;
  wire [0:0] fork84_outs_0;
  wire  fork84_outs_0_valid;
  wire  fork84_outs_0_ready;
  wire [0:0] fork84_outs_1;
  wire  fork84_outs_1_valid;
  wire  fork84_outs_1_ready;
  wire [0:0] fork84_outs_2;
  wire  fork84_outs_2_valid;
  wire  fork84_outs_2_ready;
  wire [0:0] fork84_outs_3;
  wire  fork84_outs_3_valid;
  wire  fork84_outs_3_ready;
  wire [0:0] fork84_outs_4;
  wire  fork84_outs_4_valid;
  wire  fork84_outs_4_ready;
  wire [0:0] fork84_outs_5;
  wire  fork84_outs_5_valid;
  wire  fork84_outs_5_ready;
  wire [0:0] fork84_outs_6;
  wire  fork84_outs_6_valid;
  wire  fork84_outs_6_ready;
  wire [0:0] fork84_outs_7;
  wire  fork84_outs_7_valid;
  wire  fork84_outs_7_ready;
  wire [0:0] fork84_outs_8;
  wire  fork84_outs_8_valid;
  wire  fork84_outs_8_ready;
  wire [36:0] cond_br275_trueOut;
  wire  cond_br275_trueOut_valid;
  wire  cond_br275_trueOut_ready;
  wire [36:0] cond_br275_falseOut;
  wire  cond_br275_falseOut_valid;
  wire  cond_br275_falseOut_ready;
  wire [26:0] cond_br276_trueOut;
  wire  cond_br276_trueOut_valid;
  wire  cond_br276_trueOut_ready;
  wire [26:0] cond_br276_falseOut;
  wire  cond_br276_falseOut_valid;
  wire  cond_br276_falseOut_ready;
  wire [32:0] extsi226_outs;
  wire  extsi226_outs_valid;
  wire  extsi226_outs_ready;
  wire [26:0] cond_br277_trueOut;
  wire  cond_br277_trueOut_valid;
  wire  cond_br277_trueOut_ready;
  wire [26:0] cond_br277_falseOut;
  wire  cond_br277_falseOut_valid;
  wire  cond_br277_falseOut_ready;
  wire [17:0] cond_br278_trueOut;
  wire  cond_br278_trueOut_valid;
  wire  cond_br278_trueOut_ready;
  wire [17:0] cond_br278_falseOut;
  wire  cond_br278_falseOut_valid;
  wire  cond_br278_falseOut_ready;
  wire [21:0] extsi227_outs;
  wire  extsi227_outs_valid;
  wire  extsi227_outs_ready;
  wire [16:0] cond_br279_trueOut;
  wire  cond_br279_trueOut_valid;
  wire  cond_br279_trueOut_ready;
  wire [16:0] cond_br279_falseOut;
  wire  cond_br279_falseOut_valid;
  wire  cond_br279_falseOut_ready;
  wire [6:0] cond_br280_trueOut;
  wire  cond_br280_trueOut_valid;
  wire  cond_br280_trueOut_ready;
  wire [6:0] cond_br280_falseOut;
  wire  cond_br280_falseOut_valid;
  wire  cond_br280_falseOut_ready;
  wire [11:0] extsi228_outs;
  wire  extsi228_outs_valid;
  wire  extsi228_outs_ready;
  wire [6:0] buffer156_outs;
  wire  buffer156_outs_valid;
  wire  buffer156_outs_ready;
  wire [6:0] buffer157_outs;
  wire  buffer157_outs_valid;
  wire  buffer157_outs_ready;
  wire [6:0] cond_br281_trueOut;
  wire  cond_br281_trueOut_valid;
  wire  cond_br281_trueOut_ready;
  wire [6:0] cond_br281_falseOut;
  wire  cond_br281_falseOut_valid;
  wire  cond_br281_falseOut_ready;
  wire  cond_br282_trueOut_valid;
  wire  cond_br282_trueOut_ready;
  wire  cond_br282_falseOut_valid;
  wire  cond_br282_falseOut_ready;
  wire [4:0] cond_br283_trueOut;
  wire  cond_br283_trueOut_valid;
  wire  cond_br283_trueOut_ready;
  wire [4:0] cond_br283_falseOut;
  wire  cond_br283_falseOut_valid;
  wire  cond_br283_falseOut_ready;
  wire [4:0] buffer164_outs;
  wire  buffer164_outs_valid;
  wire  buffer164_outs_ready;
  wire [4:0] buffer165_outs;
  wire  buffer165_outs_valid;
  wire  buffer165_outs_ready;
  wire [4:0] fork85_outs_0;
  wire  fork85_outs_0_valid;
  wire  fork85_outs_0_ready;
  wire [4:0] fork85_outs_1;
  wire  fork85_outs_1_valid;
  wire  fork85_outs_1_ready;
  wire [5:0] extsi229_outs;
  wire  extsi229_outs_valid;
  wire  extsi229_outs_ready;
  wire  buffer166_outs_valid;
  wire  buffer166_outs_ready;
  wire  buffer167_outs_valid;
  wire  buffer167_outs_ready;
  wire  fork86_outs_0_valid;
  wire  fork86_outs_0_ready;
  wire  fork86_outs_1_valid;
  wire  fork86_outs_1_ready;
  wire  fork86_outs_2_valid;
  wire  fork86_outs_2_ready;
  wire  fork86_outs_3_valid;
  wire  fork86_outs_3_ready;
  wire  fork86_outs_4_valid;
  wire  fork86_outs_4_ready;
  wire  fork86_outs_5_valid;
  wire  fork86_outs_5_ready;
  wire  fork86_outs_6_valid;
  wire  fork86_outs_6_ready;
  wire [36:0] constant419_outs;
  wire  constant419_outs_valid;
  wire  constant419_outs_ready;
  wire [26:0] constant556_outs;
  wire  constant556_outs_valid;
  wire  constant556_outs_ready;
  wire [26:0] constant421_outs;
  wire  constant421_outs_valid;
  wire  constant421_outs_ready;
  wire [17:0] constant557_outs;
  wire  constant557_outs_valid;
  wire  constant557_outs_ready;
  wire [16:0] constant423_outs;
  wire  constant423_outs_valid;
  wire  constant423_outs_ready;
  wire [5:0] constant558_outs;
  wire  constant558_outs_valid;
  wire  constant558_outs_ready;
  wire  source29_outs_valid;
  wire  source29_outs_ready;
  wire [5:0] constant559_outs;
  wire  constant559_outs_valid;
  wire  constant559_outs_ready;
  wire [0:0] cmpi28_result;
  wire  cmpi28_result_valid;
  wire  cmpi28_result_ready;
  wire [0:0] fork87_outs_0;
  wire  fork87_outs_0_valid;
  wire  fork87_outs_0_ready;
  wire [0:0] fork87_outs_1;
  wire  fork87_outs_1_valid;
  wire  fork87_outs_1_ready;
  wire [0:0] fork87_outs_2;
  wire  fork87_outs_2_valid;
  wire  fork87_outs_2_ready;
  wire [0:0] fork87_outs_3;
  wire  fork87_outs_3_valid;
  wire  fork87_outs_3_ready;
  wire [0:0] fork87_outs_4;
  wire  fork87_outs_4_valid;
  wire  fork87_outs_4_ready;
  wire [0:0] fork87_outs_5;
  wire  fork87_outs_5_valid;
  wire  fork87_outs_5_ready;
  wire [0:0] fork87_outs_6;
  wire  fork87_outs_6_valid;
  wire  fork87_outs_6_ready;
  wire [0:0] fork87_outs_7;
  wire  fork87_outs_7_valid;
  wire  fork87_outs_7_ready;
  wire [0:0] fork87_outs_8;
  wire  fork87_outs_8_valid;
  wire  fork87_outs_8_ready;
  wire [36:0] cond_br284_trueOut;
  wire  cond_br284_trueOut_valid;
  wire  cond_br284_trueOut_ready;
  wire [36:0] cond_br284_falseOut;
  wire  cond_br284_falseOut_valid;
  wire  cond_br284_falseOut_ready;
  wire [26:0] cond_br285_trueOut;
  wire  cond_br285_trueOut_valid;
  wire  cond_br285_trueOut_ready;
  wire [26:0] cond_br285_falseOut;
  wire  cond_br285_falseOut_valid;
  wire  cond_br285_falseOut_ready;
  wire [32:0] extsi230_outs;
  wire  extsi230_outs_valid;
  wire  extsi230_outs_ready;
  wire [26:0] cond_br286_trueOut;
  wire  cond_br286_trueOut_valid;
  wire  cond_br286_trueOut_ready;
  wire [26:0] cond_br286_falseOut;
  wire  cond_br286_falseOut_valid;
  wire  cond_br286_falseOut_ready;
  wire [17:0] cond_br287_trueOut;
  wire  cond_br287_trueOut_valid;
  wire  cond_br287_trueOut_ready;
  wire [17:0] cond_br287_falseOut;
  wire  cond_br287_falseOut_valid;
  wire  cond_br287_falseOut_ready;
  wire [21:0] extsi231_outs;
  wire  extsi231_outs_valid;
  wire  extsi231_outs_ready;
  wire [16:0] cond_br288_trueOut;
  wire  cond_br288_trueOut_valid;
  wire  cond_br288_trueOut_ready;
  wire [16:0] cond_br288_falseOut;
  wire  cond_br288_falseOut_valid;
  wire  cond_br288_falseOut_ready;
  wire [5:0] cond_br289_trueOut;
  wire  cond_br289_trueOut_valid;
  wire  cond_br289_trueOut_ready;
  wire [5:0] cond_br289_falseOut;
  wire  cond_br289_falseOut_valid;
  wire  cond_br289_falseOut_ready;
  wire [11:0] extsi232_outs;
  wire  extsi232_outs_valid;
  wire  extsi232_outs_ready;
  wire [6:0] buffer162_outs;
  wire  buffer162_outs_valid;
  wire  buffer162_outs_ready;
  wire [6:0] buffer163_outs;
  wire  buffer163_outs_valid;
  wire  buffer163_outs_ready;
  wire [6:0] cond_br290_trueOut;
  wire  cond_br290_trueOut_valid;
  wire  cond_br290_trueOut_ready;
  wire [6:0] cond_br290_falseOut;
  wire  cond_br290_falseOut_valid;
  wire  cond_br290_falseOut_ready;
  wire  cond_br291_trueOut_valid;
  wire  cond_br291_trueOut_ready;
  wire  cond_br291_falseOut_valid;
  wire  cond_br291_falseOut_ready;
  wire [4:0] cond_br292_trueOut;
  wire  cond_br292_trueOut_valid;
  wire  cond_br292_trueOut_ready;
  wire [4:0] cond_br292_falseOut;
  wire  cond_br292_falseOut_valid;
  wire  cond_br292_falseOut_ready;
  wire [4:0] buffer170_outs;
  wire  buffer170_outs_valid;
  wire  buffer170_outs_ready;
  wire [4:0] buffer171_outs;
  wire  buffer171_outs_valid;
  wire  buffer171_outs_ready;
  wire [4:0] fork88_outs_0;
  wire  fork88_outs_0_valid;
  wire  fork88_outs_0_ready;
  wire [4:0] fork88_outs_1;
  wire  fork88_outs_1_valid;
  wire  fork88_outs_1_ready;
  wire [5:0] extsi233_outs;
  wire  extsi233_outs_valid;
  wire  extsi233_outs_ready;
  wire  buffer172_outs_valid;
  wire  buffer172_outs_ready;
  wire  buffer173_outs_valid;
  wire  buffer173_outs_ready;
  wire  fork89_outs_0_valid;
  wire  fork89_outs_0_ready;
  wire  fork89_outs_1_valid;
  wire  fork89_outs_1_ready;
  wire  fork89_outs_2_valid;
  wire  fork89_outs_2_ready;
  wire  fork89_outs_3_valid;
  wire  fork89_outs_3_ready;
  wire  fork89_outs_4_valid;
  wire  fork89_outs_4_ready;
  wire  fork89_outs_5_valid;
  wire  fork89_outs_5_ready;
  wire  fork89_outs_6_valid;
  wire  fork89_outs_6_ready;
  wire [36:0] constant426_outs;
  wire  constant426_outs_valid;
  wire  constant426_outs_ready;
  wire [26:0] constant560_outs;
  wire  constant560_outs_valid;
  wire  constant560_outs_ready;
  wire [26:0] constant428_outs;
  wire  constant428_outs_valid;
  wire  constant428_outs_ready;
  wire [16:0] constant561_outs;
  wire  constant561_outs_valid;
  wire  constant561_outs_ready;
  wire [16:0] constant430_outs;
  wire  constant430_outs_valid;
  wire  constant430_outs_ready;
  wire [5:0] constant562_outs;
  wire  constant562_outs_valid;
  wire  constant562_outs_ready;
  wire  source30_outs_valid;
  wire  source30_outs_ready;
  wire [5:0] constant563_outs;
  wire  constant563_outs_valid;
  wire  constant563_outs_ready;
  wire [0:0] cmpi29_result;
  wire  cmpi29_result_valid;
  wire  cmpi29_result_ready;
  wire [0:0] fork90_outs_0;
  wire  fork90_outs_0_valid;
  wire  fork90_outs_0_ready;
  wire [0:0] fork90_outs_1;
  wire  fork90_outs_1_valid;
  wire  fork90_outs_1_ready;
  wire [0:0] fork90_outs_2;
  wire  fork90_outs_2_valid;
  wire  fork90_outs_2_ready;
  wire [0:0] fork90_outs_3;
  wire  fork90_outs_3_valid;
  wire  fork90_outs_3_ready;
  wire [0:0] fork90_outs_4;
  wire  fork90_outs_4_valid;
  wire  fork90_outs_4_ready;
  wire [0:0] fork90_outs_5;
  wire  fork90_outs_5_valid;
  wire  fork90_outs_5_ready;
  wire [0:0] fork90_outs_6;
  wire  fork90_outs_6_valid;
  wire  fork90_outs_6_ready;
  wire [0:0] fork90_outs_7;
  wire  fork90_outs_7_valid;
  wire  fork90_outs_7_ready;
  wire [0:0] fork90_outs_8;
  wire  fork90_outs_8_valid;
  wire  fork90_outs_8_ready;
  wire [36:0] cond_br293_trueOut;
  wire  cond_br293_trueOut_valid;
  wire  cond_br293_trueOut_ready;
  wire [36:0] cond_br293_falseOut;
  wire  cond_br293_falseOut_valid;
  wire  cond_br293_falseOut_ready;
  wire [26:0] cond_br294_trueOut;
  wire  cond_br294_trueOut_valid;
  wire  cond_br294_trueOut_ready;
  wire [26:0] cond_br294_falseOut;
  wire  cond_br294_falseOut_valid;
  wire  cond_br294_falseOut_ready;
  wire [32:0] extsi234_outs;
  wire  extsi234_outs_valid;
  wire  extsi234_outs_ready;
  wire [26:0] cond_br295_trueOut;
  wire  cond_br295_trueOut_valid;
  wire  cond_br295_trueOut_ready;
  wire [26:0] cond_br295_falseOut;
  wire  cond_br295_falseOut_valid;
  wire  cond_br295_falseOut_ready;
  wire [16:0] cond_br296_trueOut;
  wire  cond_br296_trueOut_valid;
  wire  cond_br296_trueOut_ready;
  wire [16:0] cond_br296_falseOut;
  wire  cond_br296_falseOut_valid;
  wire  cond_br296_falseOut_ready;
  wire [21:0] extsi235_outs;
  wire  extsi235_outs_valid;
  wire  extsi235_outs_ready;
  wire [16:0] cond_br297_trueOut;
  wire  cond_br297_trueOut_valid;
  wire  cond_br297_trueOut_ready;
  wire [16:0] cond_br297_falseOut;
  wire  cond_br297_falseOut_valid;
  wire  cond_br297_falseOut_ready;
  wire [5:0] cond_br298_trueOut;
  wire  cond_br298_trueOut_valid;
  wire  cond_br298_trueOut_ready;
  wire [5:0] cond_br298_falseOut;
  wire  cond_br298_falseOut_valid;
  wire  cond_br298_falseOut_ready;
  wire [11:0] extsi236_outs;
  wire  extsi236_outs_valid;
  wire  extsi236_outs_ready;
  wire [6:0] buffer168_outs;
  wire  buffer168_outs_valid;
  wire  buffer168_outs_ready;
  wire [6:0] buffer169_outs;
  wire  buffer169_outs_valid;
  wire  buffer169_outs_ready;
  wire [6:0] cond_br299_trueOut;
  wire  cond_br299_trueOut_valid;
  wire  cond_br299_trueOut_ready;
  wire [6:0] cond_br299_falseOut;
  wire  cond_br299_falseOut_valid;
  wire  cond_br299_falseOut_ready;
  wire  cond_br300_trueOut_valid;
  wire  cond_br300_trueOut_ready;
  wire  cond_br300_falseOut_valid;
  wire  cond_br300_falseOut_ready;
  wire [4:0] cond_br301_trueOut;
  wire  cond_br301_trueOut_valid;
  wire  cond_br301_trueOut_ready;
  wire [4:0] cond_br301_falseOut;
  wire  cond_br301_falseOut_valid;
  wire  cond_br301_falseOut_ready;
  wire [4:0] buffer176_outs;
  wire  buffer176_outs_valid;
  wire  buffer176_outs_ready;
  wire [4:0] buffer177_outs;
  wire  buffer177_outs_valid;
  wire  buffer177_outs_ready;
  wire [4:0] fork91_outs_0;
  wire  fork91_outs_0_valid;
  wire  fork91_outs_0_ready;
  wire [4:0] fork91_outs_1;
  wire  fork91_outs_1_valid;
  wire  fork91_outs_1_ready;
  wire [5:0] extsi237_outs;
  wire  extsi237_outs_valid;
  wire  extsi237_outs_ready;
  wire  buffer178_outs_valid;
  wire  buffer178_outs_ready;
  wire  buffer179_outs_valid;
  wire  buffer179_outs_ready;
  wire  fork92_outs_0_valid;
  wire  fork92_outs_0_ready;
  wire  fork92_outs_1_valid;
  wire  fork92_outs_1_ready;
  wire  fork92_outs_2_valid;
  wire  fork92_outs_2_ready;
  wire  fork92_outs_3_valid;
  wire  fork92_outs_3_ready;
  wire  fork92_outs_4_valid;
  wire  fork92_outs_4_ready;
  wire  fork92_outs_5_valid;
  wire  fork92_outs_5_ready;
  wire  fork92_outs_6_valid;
  wire  fork92_outs_6_ready;
  wire [36:0] constant433_outs;
  wire  constant433_outs_valid;
  wire  constant433_outs_ready;
  wire [26:0] constant564_outs;
  wire  constant564_outs_valid;
  wire  constant564_outs_ready;
  wire [26:0] constant435_outs;
  wire  constant435_outs_valid;
  wire  constant435_outs_ready;
  wire [16:0] constant565_outs;
  wire  constant565_outs_valid;
  wire  constant565_outs_ready;
  wire [16:0] constant437_outs;
  wire  constant437_outs_valid;
  wire  constant437_outs_ready;
  wire [5:0] constant566_outs;
  wire  constant566_outs_valid;
  wire  constant566_outs_ready;
  wire  source31_outs_valid;
  wire  source31_outs_ready;
  wire [5:0] constant567_outs;
  wire  constant567_outs_valid;
  wire  constant567_outs_ready;
  wire [0:0] cmpi30_result;
  wire  cmpi30_result_valid;
  wire  cmpi30_result_ready;
  wire [0:0] fork93_outs_0;
  wire  fork93_outs_0_valid;
  wire  fork93_outs_0_ready;
  wire [0:0] fork93_outs_1;
  wire  fork93_outs_1_valid;
  wire  fork93_outs_1_ready;
  wire [0:0] fork93_outs_2;
  wire  fork93_outs_2_valid;
  wire  fork93_outs_2_ready;
  wire [0:0] fork93_outs_3;
  wire  fork93_outs_3_valid;
  wire  fork93_outs_3_ready;
  wire [0:0] fork93_outs_4;
  wire  fork93_outs_4_valid;
  wire  fork93_outs_4_ready;
  wire [0:0] fork93_outs_5;
  wire  fork93_outs_5_valid;
  wire  fork93_outs_5_ready;
  wire [0:0] fork93_outs_6;
  wire  fork93_outs_6_valid;
  wire  fork93_outs_6_ready;
  wire [0:0] fork93_outs_7;
  wire  fork93_outs_7_valid;
  wire  fork93_outs_7_ready;
  wire [0:0] fork93_outs_8;
  wire  fork93_outs_8_valid;
  wire  fork93_outs_8_ready;
  wire [36:0] cond_br302_trueOut;
  wire  cond_br302_trueOut_valid;
  wire  cond_br302_trueOut_ready;
  wire [36:0] cond_br302_falseOut;
  wire  cond_br302_falseOut_valid;
  wire  cond_br302_falseOut_ready;
  wire [26:0] cond_br303_trueOut;
  wire  cond_br303_trueOut_valid;
  wire  cond_br303_trueOut_ready;
  wire [26:0] cond_br303_falseOut;
  wire  cond_br303_falseOut_valid;
  wire  cond_br303_falseOut_ready;
  wire [32:0] extsi238_outs;
  wire  extsi238_outs_valid;
  wire  extsi238_outs_ready;
  wire [26:0] cond_br304_trueOut;
  wire  cond_br304_trueOut_valid;
  wire  cond_br304_trueOut_ready;
  wire [26:0] cond_br304_falseOut;
  wire  cond_br304_falseOut_valid;
  wire  cond_br304_falseOut_ready;
  wire [16:0] cond_br305_trueOut;
  wire  cond_br305_trueOut_valid;
  wire  cond_br305_trueOut_ready;
  wire [16:0] cond_br305_falseOut;
  wire  cond_br305_falseOut_valid;
  wire  cond_br305_falseOut_ready;
  wire [21:0] extsi239_outs;
  wire  extsi239_outs_valid;
  wire  extsi239_outs_ready;
  wire [16:0] cond_br306_trueOut;
  wire  cond_br306_trueOut_valid;
  wire  cond_br306_trueOut_ready;
  wire [16:0] cond_br306_falseOut;
  wire  cond_br306_falseOut_valid;
  wire  cond_br306_falseOut_ready;
  wire [5:0] cond_br307_trueOut;
  wire  cond_br307_trueOut_valid;
  wire  cond_br307_trueOut_ready;
  wire [5:0] cond_br307_falseOut;
  wire  cond_br307_falseOut_valid;
  wire  cond_br307_falseOut_ready;
  wire [11:0] extsi240_outs;
  wire  extsi240_outs_valid;
  wire  extsi240_outs_ready;
  wire [6:0] buffer174_outs;
  wire  buffer174_outs_valid;
  wire  buffer174_outs_ready;
  wire [6:0] buffer175_outs;
  wire  buffer175_outs_valid;
  wire  buffer175_outs_ready;
  wire [6:0] cond_br308_trueOut;
  wire  cond_br308_trueOut_valid;
  wire  cond_br308_trueOut_ready;
  wire [6:0] cond_br308_falseOut;
  wire  cond_br308_falseOut_valid;
  wire  cond_br308_falseOut_ready;
  wire  cond_br309_trueOut_valid;
  wire  cond_br309_trueOut_ready;
  wire  cond_br309_falseOut_valid;
  wire  cond_br309_falseOut_ready;
  wire [4:0] cond_br310_trueOut;
  wire  cond_br310_trueOut_valid;
  wire  cond_br310_trueOut_ready;
  wire [4:0] cond_br310_falseOut;
  wire  cond_br310_falseOut_valid;
  wire  cond_br310_falseOut_ready;
  wire [4:0] buffer182_outs;
  wire  buffer182_outs_valid;
  wire  buffer182_outs_ready;
  wire [4:0] buffer183_outs;
  wire  buffer183_outs_valid;
  wire  buffer183_outs_ready;
  wire [5:0] extsi241_outs;
  wire  extsi241_outs_valid;
  wire  extsi241_outs_ready;
  wire  buffer184_outs_valid;
  wire  buffer184_outs_ready;
  wire  buffer185_outs_valid;
  wire  buffer185_outs_ready;
  wire  fork94_outs_0_valid;
  wire  fork94_outs_0_ready;
  wire  fork94_outs_1_valid;
  wire  fork94_outs_1_ready;
  wire  fork94_outs_2_valid;
  wire  fork94_outs_2_ready;
  wire  fork94_outs_3_valid;
  wire  fork94_outs_3_ready;
  wire  fork94_outs_4_valid;
  wire  fork94_outs_4_ready;
  wire  fork94_outs_5_valid;
  wire  fork94_outs_5_ready;
  wire  fork94_outs_6_valid;
  wire  fork94_outs_6_ready;
  wire  fork94_outs_7_valid;
  wire  fork94_outs_7_ready;
  wire  fork94_outs_8_valid;
  wire  fork94_outs_8_ready;
  wire  fork94_outs_9_valid;
  wire  fork94_outs_9_ready;
  wire  fork94_outs_10_valid;
  wire  fork94_outs_10_ready;
  wire  fork94_outs_11_valid;
  wire  fork94_outs_11_ready;
  wire  fork94_outs_12_valid;
  wire  fork94_outs_12_ready;
  wire [32:0] constant568_outs;
  wire  constant568_outs_valid;
  wire  constant568_outs_ready;
  wire [32:0] constant441_outs;
  wire  constant441_outs_valid;
  wire  constant441_outs_ready;
  wire [26:0] constant442_outs;
  wire  constant442_outs_valid;
  wire  constant442_outs_ready;
  wire [21:0] constant443_outs;
  wire  constant443_outs_valid;
  wire  constant443_outs_ready;
  wire [14:0] constant569_outs;
  wire  constant569_outs_valid;
  wire  constant569_outs_ready;
  wire [11:0] constant445_outs;
  wire  constant445_outs_valid;
  wire  constant445_outs_ready;
  wire [36:0] constant446_outs;
  wire  constant446_outs_valid;
  wire  constant446_outs_ready;
  wire [25:0] constant570_outs;
  wire  constant570_outs_valid;
  wire  constant570_outs_ready;
  wire [26:0] constant448_outs;
  wire  constant448_outs_valid;
  wire  constant448_outs_ready;
  wire [16:0] constant571_outs;
  wire  constant571_outs_valid;
  wire  constant571_outs_ready;
  wire [16:0] constant450_outs;
  wire  constant450_outs_valid;
  wire  constant450_outs_ready;
  wire [5:0] constant572_outs;
  wire  constant572_outs_valid;
  wire  constant572_outs_ready;
  wire  source32_outs_valid;
  wire  source32_outs_ready;
  wire [5:0] constant573_outs;
  wire  constant573_outs_valid;
  wire  constant573_outs_ready;
  wire [0:0] cmpi31_result;
  wire  cmpi31_result_valid;
  wire  cmpi31_result_ready;
  wire [0:0] fork95_outs_0;
  wire  fork95_outs_0_valid;
  wire  fork95_outs_0_ready;
  wire [0:0] fork95_outs_1;
  wire  fork95_outs_1_valid;
  wire  fork95_outs_1_ready;
  wire [0:0] fork95_outs_2;
  wire  fork95_outs_2_valid;
  wire  fork95_outs_2_ready;
  wire [0:0] fork95_outs_3;
  wire  fork95_outs_3_valid;
  wire  fork95_outs_3_ready;
  wire [0:0] fork95_outs_4;
  wire  fork95_outs_4_valid;
  wire  fork95_outs_4_ready;
  wire [0:0] fork95_outs_5;
  wire  fork95_outs_5_valid;
  wire  fork95_outs_5_ready;
  wire [0:0] fork95_outs_6;
  wire  fork95_outs_6_valid;
  wire  fork95_outs_6_ready;
  wire [0:0] fork95_outs_7;
  wire  fork95_outs_7_valid;
  wire  fork95_outs_7_ready;
  wire [0:0] fork95_outs_8;
  wire  fork95_outs_8_valid;
  wire  fork95_outs_8_ready;
  wire [0:0] fork95_outs_9;
  wire  fork95_outs_9_valid;
  wire  fork95_outs_9_ready;
  wire [0:0] fork95_outs_10;
  wire  fork95_outs_10_valid;
  wire  fork95_outs_10_ready;
  wire [0:0] fork95_outs_11;
  wire  fork95_outs_11_valid;
  wire  fork95_outs_11_ready;
  wire [0:0] fork95_outs_12;
  wire  fork95_outs_12_valid;
  wire  fork95_outs_12_ready;
  wire [0:0] fork95_outs_13;
  wire  fork95_outs_13_valid;
  wire  fork95_outs_13_ready;
  wire [36:0] cond_br311_trueOut;
  wire  cond_br311_trueOut_valid;
  wire  cond_br311_trueOut_ready;
  wire [36:0] cond_br311_falseOut;
  wire  cond_br311_falseOut_valid;
  wire  cond_br311_falseOut_ready;
  wire [25:0] cond_br312_trueOut;
  wire  cond_br312_trueOut_valid;
  wire  cond_br312_trueOut_ready;
  wire [25:0] cond_br312_falseOut;
  wire  cond_br312_falseOut_valid;
  wire  cond_br312_falseOut_ready;
  wire [32:0] extsi242_outs;
  wire  extsi242_outs_valid;
  wire  extsi242_outs_ready;
  wire [26:0] cond_br313_trueOut;
  wire  cond_br313_trueOut_valid;
  wire  cond_br313_trueOut_ready;
  wire [26:0] cond_br313_falseOut;
  wire  cond_br313_falseOut_valid;
  wire  cond_br313_falseOut_ready;
  wire [16:0] cond_br314_trueOut;
  wire  cond_br314_trueOut_valid;
  wire  cond_br314_trueOut_ready;
  wire [16:0] cond_br314_falseOut;
  wire  cond_br314_falseOut_valid;
  wire  cond_br314_falseOut_ready;
  wire [21:0] extsi243_outs;
  wire  extsi243_outs_valid;
  wire  extsi243_outs_ready;
  wire [16:0] cond_br315_trueOut;
  wire  cond_br315_trueOut_valid;
  wire  cond_br315_trueOut_ready;
  wire [16:0] cond_br315_falseOut;
  wire  cond_br315_falseOut_valid;
  wire  cond_br315_falseOut_ready;
  wire [5:0] cond_br316_trueOut;
  wire  cond_br316_trueOut_valid;
  wire  cond_br316_trueOut_ready;
  wire [5:0] cond_br316_falseOut;
  wire  cond_br316_falseOut_valid;
  wire  cond_br316_falseOut_ready;
  wire [11:0] extsi244_outs;
  wire  extsi244_outs_valid;
  wire  extsi244_outs_ready;
  wire [6:0] buffer180_outs;
  wire  buffer180_outs_valid;
  wire  buffer180_outs_ready;
  wire [6:0] buffer181_outs;
  wire  buffer181_outs_valid;
  wire  buffer181_outs_ready;
  wire [6:0] cond_br317_trueOut;
  wire  cond_br317_trueOut_valid;
  wire  cond_br317_trueOut_ready;
  wire [6:0] cond_br317_falseOut;
  wire  cond_br317_falseOut_valid;
  wire  cond_br317_falseOut_ready;
  wire [6:0] fork96_outs_0;
  wire  fork96_outs_0_valid;
  wire  fork96_outs_0_ready;
  wire [6:0] fork96_outs_1;
  wire  fork96_outs_1_valid;
  wire  fork96_outs_1_ready;
  wire  cond_br318_trueOut_valid;
  wire  cond_br318_trueOut_ready;
  wire  cond_br318_falseOut_valid;
  wire  cond_br318_falseOut_ready;
  wire  fork97_outs_0_valid;
  wire  fork97_outs_0_ready;
  wire  fork97_outs_1_valid;
  wire  fork97_outs_1_ready;
  wire [32:0] cond_br319_trueOut;
  wire  cond_br319_trueOut_valid;
  wire  cond_br319_trueOut_ready;
  wire [32:0] cond_br319_falseOut;
  wire  cond_br319_falseOut_valid;
  wire  cond_br319_falseOut_ready;
  wire [36:0] extsi245_outs;
  wire  extsi245_outs_valid;
  wire  extsi245_outs_ready;
  wire [32:0] cond_br320_trueOut;
  wire  cond_br320_trueOut_valid;
  wire  cond_br320_trueOut_ready;
  wire [32:0] cond_br320_falseOut;
  wire  cond_br320_falseOut_valid;
  wire  cond_br320_falseOut_ready;
  wire [26:0] cond_br321_trueOut;
  wire  cond_br321_trueOut_valid;
  wire  cond_br321_trueOut_ready;
  wire [26:0] cond_br321_falseOut;
  wire  cond_br321_falseOut_valid;
  wire  cond_br321_falseOut_ready;
  wire [21:0] cond_br322_trueOut;
  wire  cond_br322_trueOut_valid;
  wire  cond_br322_trueOut_ready;
  wire [21:0] cond_br322_falseOut;
  wire  cond_br322_falseOut_valid;
  wire  cond_br322_falseOut_ready;
  wire [14:0] cond_br323_trueOut;
  wire  cond_br323_trueOut_valid;
  wire  cond_br323_trueOut_ready;
  wire [14:0] cond_br323_falseOut;
  wire  cond_br323_falseOut_valid;
  wire  cond_br323_falseOut_ready;
  wire [16:0] extsi246_outs;
  wire  extsi246_outs_valid;
  wire  extsi246_outs_ready;
  wire [11:0] cond_br324_trueOut;
  wire  cond_br324_trueOut_valid;
  wire  cond_br324_trueOut_ready;
  wire [11:0] cond_br324_falseOut;
  wire  cond_br324_falseOut_valid;
  wire  cond_br324_falseOut_ready;
  wire [36:0] mux0_outs;
  wire  mux0_outs_valid;
  wire  mux0_outs_ready;
  wire [32:0] mux1_outs;
  wire  mux1_outs_valid;
  wire  mux1_outs_ready;
  wire [26:0] mux2_outs;
  wire  mux2_outs_valid;
  wire  mux2_outs_ready;
  wire [21:0] mux3_outs;
  wire  mux3_outs_valid;
  wire  mux3_outs_ready;
  wire [16:0] mux4_outs;
  wire  mux4_outs_valid;
  wire  mux4_outs_ready;
  wire [11:0] mux5_outs;
  wire  mux5_outs_valid;
  wire  mux5_outs_ready;
  wire [6:0] mux6_outs;
  wire  mux6_outs_valid;
  wire  mux6_outs_ready;
  wire [6:0] buffer198_outs;
  wire  buffer198_outs_valid;
  wire  buffer198_outs_ready;
  wire [6:0] buffer199_outs;
  wire  buffer199_outs_valid;
  wire  buffer199_outs_ready;
  wire [6:0] fork98_outs_0;
  wire  fork98_outs_0_valid;
  wire  fork98_outs_0_ready;
  wire [6:0] fork98_outs_1;
  wire  fork98_outs_1_valid;
  wire  fork98_outs_1_ready;
  wire [6:0] fork98_outs_2;
  wire  fork98_outs_2_valid;
  wire  fork98_outs_2_ready;
  wire [6:0] fork98_outs_3;
  wire  fork98_outs_3_valid;
  wire  fork98_outs_3_ready;
  wire [6:0] fork98_outs_4;
  wire  fork98_outs_4_valid;
  wire  fork98_outs_4_ready;
  wire  control_merge31_outs_valid;
  wire  control_merge31_outs_ready;
  wire [5:0] control_merge31_index;
  wire  control_merge31_index_valid;
  wire  control_merge31_index_ready;
  wire [5:0] fork99_outs_0;
  wire  fork99_outs_0_valid;
  wire  fork99_outs_0_ready;
  wire [5:0] fork99_outs_1;
  wire  fork99_outs_1_valid;
  wire  fork99_outs_1_ready;
  wire [5:0] fork99_outs_2;
  wire  fork99_outs_2_valid;
  wire  fork99_outs_2_ready;
  wire [5:0] fork99_outs_3;
  wire  fork99_outs_3_valid;
  wire  fork99_outs_3_ready;
  wire [5:0] fork99_outs_4;
  wire  fork99_outs_4_valid;
  wire  fork99_outs_4_ready;
  wire [5:0] fork99_outs_5;
  wire  fork99_outs_5_valid;
  wire  fork99_outs_5_ready;
  wire [5:0] fork99_outs_6;
  wire  fork99_outs_6_valid;
  wire  fork99_outs_6_ready;
  wire  buffer200_outs_valid;
  wire  buffer200_outs_ready;
  wire  buffer201_outs_valid;
  wire  buffer201_outs_ready;
  wire  source33_outs_valid;
  wire  source33_outs_ready;
  wire [1:0] constant574_outs;
  wire  constant574_outs_valid;
  wire  constant574_outs_ready;
  wire [1:0] fork100_outs_0;
  wire  fork100_outs_0_valid;
  wire  fork100_outs_0_ready;
  wire [1:0] fork100_outs_1;
  wire  fork100_outs_1_valid;
  wire  fork100_outs_1_ready;
  wire [1:0] fork100_outs_2;
  wire  fork100_outs_2_valid;
  wire  fork100_outs_2_ready;
  wire [1:0] fork100_outs_3;
  wire  fork100_outs_3_valid;
  wire  fork100_outs_3_ready;
  wire [1:0] fork100_outs_4;
  wire  fork100_outs_4_valid;
  wire  fork100_outs_4_ready;
  wire [38:0] extsi135_outs;
  wire  extsi135_outs_valid;
  wire  extsi135_outs_ready;
  wire [34:0] extsi136_outs;
  wire  extsi136_outs_valid;
  wire  extsi136_outs_ready;
  wire [28:0] extsi137_outs;
  wire  extsi137_outs_valid;
  wire  extsi137_outs_ready;
  wire [23:0] extsi138_outs;
  wire  extsi138_outs_valid;
  wire  extsi138_outs_ready;
  wire [18:0] extsi139_outs;
  wire  extsi139_outs_valid;
  wire  extsi139_outs_ready;
  wire  source38_outs_valid;
  wire  source38_outs_ready;
  wire [3:0] constant575_outs;
  wire  constant575_outs_valid;
  wire  constant575_outs_ready;
  wire [11:0] extui0_outs;
  wire  extui0_outs_valid;
  wire  extui0_outs_ready;
  wire [5:0] trunci1_outs;
  wire  trunci1_outs_valid;
  wire  trunci1_outs_ready;
  wire [11:0] buffer196_outs;
  wire  buffer196_outs_valid;
  wire  buffer196_outs_ready;
  wire [11:0] buffer197_outs;
  wire  buffer197_outs_valid;
  wire  buffer197_outs_ready;
  wire [17:0] extsi0_outs;
  wire  extsi0_outs_valid;
  wire  extsi0_outs_ready;
  wire [17:0] extsi1_outs;
  wire  extsi1_outs_valid;
  wire  extsi1_outs_ready;
  wire [17:0] muli0_result;
  wire  muli0_result_valid;
  wire  muli0_result_ready;
  wire [16:0] buffer194_outs;
  wire  buffer194_outs_valid;
  wire  buffer194_outs_ready;
  wire [16:0] buffer195_outs;
  wire  buffer195_outs_valid;
  wire  buffer195_outs_ready;
  wire [18:0] extsi3_outs;
  wire  extsi3_outs_valid;
  wire  extsi3_outs_ready;
  wire [18:0] shli0_result;
  wire  shli0_result_valid;
  wire  shli0_result_ready;
  wire [17:0] trunci14_outs;
  wire  trunci14_outs_valid;
  wire  trunci14_outs_ready;
  wire [17:0] addi0_result;
  wire  addi0_result_valid;
  wire  addi0_result_ready;
  wire [24:0] extsi4_outs;
  wire  extsi4_outs_valid;
  wire  extsi4_outs_ready;
  wire [24:0] extsi5_outs;
  wire  extsi5_outs_valid;
  wire  extsi5_outs_ready;
  wire [24:0] muli1_result;
  wire  muli1_result_valid;
  wire  muli1_result_ready;
  wire [22:0] trunci4_outs;
  wire  trunci4_outs_valid;
  wire  trunci4_outs_ready;
  wire [21:0] buffer192_outs;
  wire  buffer192_outs_valid;
  wire  buffer192_outs_ready;
  wire [21:0] buffer193_outs;
  wire  buffer193_outs_valid;
  wire  buffer193_outs_ready;
  wire [23:0] extsi7_outs;
  wire  extsi7_outs_valid;
  wire  extsi7_outs_ready;
  wire [23:0] shli1_result;
  wire  shli1_result_valid;
  wire  shli1_result_ready;
  wire [22:0] trunci15_outs;
  wire  trunci15_outs_valid;
  wire  trunci15_outs_ready;
  wire [22:0] addi1_result;
  wire  addi1_result_valid;
  wire  addi1_result_ready;
  wire [29:0] extsi8_outs;
  wire  extsi8_outs_valid;
  wire  extsi8_outs_ready;
  wire [29:0] extsi9_outs;
  wire  extsi9_outs_valid;
  wire  extsi9_outs_ready;
  wire [29:0] muli2_result;
  wire  muli2_result_valid;
  wire  muli2_result_ready;
  wire [27:0] trunci6_outs;
  wire  trunci6_outs_valid;
  wire  trunci6_outs_ready;
  wire [26:0] buffer190_outs;
  wire  buffer190_outs_valid;
  wire  buffer190_outs_ready;
  wire [26:0] buffer191_outs;
  wire  buffer191_outs_valid;
  wire  buffer191_outs_ready;
  wire [28:0] extsi11_outs;
  wire  extsi11_outs_valid;
  wire  extsi11_outs_ready;
  wire [28:0] shli2_result;
  wire  shli2_result_valid;
  wire  shli2_result_ready;
  wire [27:0] trunci16_outs;
  wire  trunci16_outs_valid;
  wire  trunci16_outs_ready;
  wire [27:0] addi2_result;
  wire  addi2_result_valid;
  wire  addi2_result_ready;
  wire [34:0] extsi12_outs;
  wire  extsi12_outs_valid;
  wire  extsi12_outs_ready;
  wire [34:0] extsi13_outs;
  wire  extsi13_outs_valid;
  wire  extsi13_outs_ready;
  wire [34:0] muli3_result;
  wire  muli3_result_valid;
  wire  muli3_result_ready;
  wire [33:0] trunci8_outs;
  wire  trunci8_outs_valid;
  wire  trunci8_outs_ready;
  wire [32:0] buffer188_outs;
  wire  buffer188_outs_valid;
  wire  buffer188_outs_ready;
  wire [32:0] buffer189_outs;
  wire  buffer189_outs_valid;
  wire  buffer189_outs_ready;
  wire [34:0] extsi15_outs;
  wire  extsi15_outs_valid;
  wire  extsi15_outs_ready;
  wire [34:0] shli3_result;
  wire  shli3_result_valid;
  wire  shli3_result_ready;
  wire [33:0] trunci17_outs;
  wire  trunci17_outs_valid;
  wire  trunci17_outs_ready;
  wire [33:0] addi3_result;
  wire  addi3_result_valid;
  wire  addi3_result_ready;
  wire [40:0] extsi16_outs;
  wire  extsi16_outs_valid;
  wire  extsi16_outs_ready;
  wire [40:0] extsi17_outs;
  wire  extsi17_outs_valid;
  wire  extsi17_outs_ready;
  wire [40:0] muli4_result;
  wire  muli4_result_valid;
  wire  muli4_result_ready;
  wire [11:0] trunci18_outs;
  wire  trunci18_outs_valid;
  wire  trunci18_outs_ready;
  wire [36:0] buffer186_outs;
  wire  buffer186_outs_valid;
  wire  buffer186_outs_ready;
  wire [36:0] buffer187_outs;
  wire  buffer187_outs_valid;
  wire  buffer187_outs_ready;
  wire [38:0] extsi19_outs;
  wire  extsi19_outs_valid;
  wire  extsi19_outs_ready;
  wire [38:0] shli4_result;
  wire  shli4_result_valid;
  wire  shli4_result_ready;
  wire [11:0] trunci19_outs;
  wire  trunci19_outs_valid;
  wire  trunci19_outs_ready;
  wire [11:0] addi4_result;
  wire  addi4_result_valid;
  wire  addi4_result_ready;
  wire [11:0] shrsi0_result;
  wire  shrsi0_result_valid;
  wire  shrsi0_result_ready;
  wire [7:0] trunci12_outs;
  wire  trunci12_outs_valid;
  wire  trunci12_outs_ready;

  assign out0 = trunci12_outs;
  assign out0_valid = trunci12_outs_valid;
  assign trunci12_outs_ready = out0_ready;
  assign end_valid = fork0_outs_6_valid;
  assign fork0_outs_6_ready = end_ready;

  fork_dataless #(.SIZE(8)) fork0(
    .ins_valid (start_valid),
    .ins_ready (start_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork0_outs_7_valid, fork0_outs_6_valid, fork0_outs_5_valid, fork0_outs_4_valid, fork0_outs_3_valid, fork0_outs_2_valid, fork0_outs_1_valid, fork0_outs_0_valid}),
    .outs_ready ({fork0_outs_7_ready, fork0_outs_6_ready, fork0_outs_5_ready, fork0_outs_4_ready, fork0_outs_3_ready, fork0_outs_2_ready, fork0_outs_1_ready, fork0_outs_0_ready})
  );

  fork_type #(.SIZE(2), .DATA_TYPE(17)) fork1(
    .ins (in0),
    .ins_valid (in0_valid),
    .ins_ready (in0_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork1_outs_1, fork1_outs_0}),
    .outs_valid ({fork1_outs_1_valid, fork1_outs_0_valid}),
    .outs_ready ({fork1_outs_1_ready, fork1_outs_0_ready})
  );

  trunci #(.INPUT_TYPE(17), .OUTPUT_TYPE(7)) trunci13(
    .ins (fork1_outs_0),
    .ins_valid (fork1_outs_0_valid),
    .ins_ready (fork1_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci13_outs),
    .outs_valid (trunci13_outs_valid),
    .outs_ready (trunci13_outs_ready)
  );

  source source0(
    .clk (clk),
    .rst (rst),
    .outs_valid (source0_outs_valid),
    .outs_ready (source0_outs_ready)
  );

  handshake_constant_0 #(.DATA_WIDTH(1)) constant459(
    .ctrl_valid (source0_outs_valid),
    .ctrl_ready (source0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant459_outs),
    .outs_valid (constant459_outs_valid),
    .outs_ready (constant459_outs_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(5)) extsi141(
    .ins (constant459_outs),
    .ins_valid (constant459_outs_valid),
    .ins_ready (constant459_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi141_outs),
    .outs_valid (extsi141_outs_valid),
    .outs_ready (extsi141_outs_ready)
  );

  handshake_constant_1 #(.DATA_WIDTH(12)) constant223(
    .ctrl_valid (fork0_outs_5_valid),
    .ctrl_ready (fork0_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant223_outs),
    .outs_valid (constant223_outs_valid),
    .outs_ready (constant223_outs_ready)
  );

  handshake_constant_2 #(.DATA_WIDTH(15)) constant460(
    .ctrl_valid (fork0_outs_1_valid),
    .ctrl_ready (fork0_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant460_outs),
    .outs_valid (constant460_outs_valid),
    .outs_ready (constant460_outs_ready)
  );

  handshake_constant_3 #(.DATA_WIDTH(22)) constant225(
    .ctrl_valid (fork0_outs_4_valid),
    .ctrl_ready (fork0_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant225_outs),
    .outs_valid (constant225_outs_valid),
    .outs_ready (constant225_outs_ready)
  );

  handshake_constant_4 #(.DATA_WIDTH(27)) constant226(
    .ctrl_valid (fork0_outs_3_valid),
    .ctrl_ready (fork0_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant226_outs),
    .outs_valid (constant226_outs_valid),
    .outs_ready (constant226_outs_ready)
  );

  handshake_constant_5 #(.DATA_WIDTH(33)) constant227(
    .ctrl_valid (fork0_outs_2_valid),
    .ctrl_ready (fork0_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant227_outs),
    .outs_valid (constant227_outs_valid),
    .outs_ready (constant227_outs_ready)
  );

  handshake_constant_6 #(.DATA_WIDTH(33)) constant461(
    .ctrl_valid (fork0_outs_0_valid),
    .ctrl_ready (fork0_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant461_outs),
    .outs_valid (constant461_outs_valid),
    .outs_ready (constant461_outs_ready)
  );

  source source1(
    .clk (clk),
    .rst (rst),
    .outs_valid (source1_outs_valid),
    .outs_ready (source1_outs_ready)
  );

  handshake_constant_7 #(.DATA_WIDTH(5)) constant462(
    .ctrl_valid (source1_outs_valid),
    .ctrl_ready (source1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant462_outs),
    .outs_valid (constant462_outs_valid),
    .outs_ready (constant462_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(17)) extsi23(
    .ins (constant462_outs),
    .ins_valid (constant462_outs_valid),
    .ins_ready (constant462_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi23_outs),
    .outs_valid (extsi23_outs_valid),
    .outs_ready (extsi23_outs_ready)
  );

  shrui #(.DATA_TYPE(17)) shrui0(
    .lhs (fork1_outs_1),
    .lhs_valid (fork1_outs_1_valid),
    .lhs_ready (fork1_outs_1_ready),
    .rhs (extsi23_outs),
    .rhs_valid (extsi23_outs_valid),
    .rhs_ready (extsi23_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shrui0_result),
    .result_valid (shrui0_result_valid),
    .result_ready (shrui0_result_ready)
  );

  trunci #(.INPUT_TYPE(17), .OUTPUT_TYPE(5)) trunci0(
    .ins (shrui0_result),
    .ins_valid (shrui0_result_valid),
    .ins_ready (shrui0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci0_outs),
    .outs_valid (trunci0_outs_valid),
    .outs_ready (trunci0_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork2(
    .ins (trunci0_outs),
    .ins_valid (trunci0_outs_valid),
    .ins_ready (trunci0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork2_outs_1, fork2_outs_0}),
    .outs_valid ({fork2_outs_1_valid, fork2_outs_0_valid}),
    .outs_ready ({fork2_outs_1_ready, fork2_outs_0_ready})
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi0(
    .lhs (fork2_outs_0),
    .lhs_valid (fork2_outs_0_valid),
    .lhs_ready (fork2_outs_0_ready),
    .rhs (extsi141_outs),
    .rhs_valid (extsi141_outs_valid),
    .rhs_ready (extsi141_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi0_result),
    .result_valid (cmpi0_result_valid),
    .result_ready (cmpi0_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork3(
    .ins (cmpi0_result),
    .ins_valid (cmpi0_result_valid),
    .ins_ready (cmpi0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork3_outs_8, fork3_outs_7, fork3_outs_6, fork3_outs_5, fork3_outs_4, fork3_outs_3, fork3_outs_2, fork3_outs_1, fork3_outs_0}),
    .outs_valid ({fork3_outs_8_valid, fork3_outs_7_valid, fork3_outs_6_valid, fork3_outs_5_valid, fork3_outs_4_valid, fork3_outs_3_valid, fork3_outs_2_valid, fork3_outs_1_valid, fork3_outs_0_valid}),
    .outs_ready ({fork3_outs_8_ready, fork3_outs_7_ready, fork3_outs_6_ready, fork3_outs_5_ready, fork3_outs_4_ready, fork3_outs_3_ready, fork3_outs_2_ready, fork3_outs_1_ready, fork3_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(33)) cond_br32(
    .condition (fork3_outs_8),
    .condition_valid (fork3_outs_8_valid),
    .condition_ready (fork3_outs_8_ready),
    .data (constant461_outs),
    .data_valid (constant461_outs_valid),
    .data_ready (constant461_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br32_trueOut),
    .trueOut_valid (cond_br32_trueOut_valid),
    .trueOut_ready (cond_br32_trueOut_ready),
    .falseOut (cond_br32_falseOut),
    .falseOut_valid (cond_br32_falseOut_valid),
    .falseOut_ready (cond_br32_falseOut_ready)
  );

  sink #(.DATA_TYPE(33)) sink0(
    .ins (cond_br32_falseOut),
    .ins_valid (cond_br32_falseOut_valid),
    .ins_ready (cond_br32_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(33), .OUTPUT_TYPE(37)) extsi142(
    .ins (cond_br32_trueOut),
    .ins_valid (cond_br32_trueOut_valid),
    .ins_ready (cond_br32_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi142_outs),
    .outs_valid (extsi142_outs_valid),
    .outs_ready (extsi142_outs_ready)
  );

  cond_br #(.DATA_TYPE(33)) cond_br33(
    .condition (fork3_outs_5),
    .condition_valid (fork3_outs_5_valid),
    .condition_ready (fork3_outs_5_ready),
    .data (constant227_outs),
    .data_valid (constant227_outs_valid),
    .data_ready (constant227_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br33_trueOut),
    .trueOut_valid (cond_br33_trueOut_valid),
    .trueOut_ready (cond_br33_trueOut_ready),
    .falseOut (cond_br33_falseOut),
    .falseOut_valid (cond_br33_falseOut_valid),
    .falseOut_ready (cond_br33_falseOut_ready)
  );

  sink #(.DATA_TYPE(33)) sink1(
    .ins (cond_br33_falseOut),
    .ins_valid (cond_br33_falseOut_valid),
    .ins_ready (cond_br33_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br34(
    .condition (fork3_outs_4),
    .condition_valid (fork3_outs_4_valid),
    .condition_ready (fork3_outs_4_ready),
    .data (constant226_outs),
    .data_valid (constant226_outs_valid),
    .data_ready (constant226_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br34_trueOut),
    .trueOut_valid (cond_br34_trueOut_valid),
    .trueOut_ready (cond_br34_trueOut_ready),
    .falseOut (cond_br34_falseOut),
    .falseOut_valid (cond_br34_falseOut_valid),
    .falseOut_ready (cond_br34_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink2(
    .ins (cond_br34_falseOut),
    .ins_valid (cond_br34_falseOut_valid),
    .ins_ready (cond_br34_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(22)) cond_br35(
    .condition (fork3_outs_3),
    .condition_valid (fork3_outs_3_valid),
    .condition_ready (fork3_outs_3_ready),
    .data (constant225_outs),
    .data_valid (constant225_outs_valid),
    .data_ready (constant225_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br35_trueOut),
    .trueOut_valid (cond_br35_trueOut_valid),
    .trueOut_ready (cond_br35_trueOut_ready),
    .falseOut (cond_br35_falseOut),
    .falseOut_valid (cond_br35_falseOut_valid),
    .falseOut_ready (cond_br35_falseOut_ready)
  );

  sink #(.DATA_TYPE(22)) sink3(
    .ins (cond_br35_falseOut),
    .ins_valid (cond_br35_falseOut_valid),
    .ins_ready (cond_br35_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(15)) cond_br36(
    .condition (fork3_outs_7),
    .condition_valid (fork3_outs_7_valid),
    .condition_ready (fork3_outs_7_ready),
    .data (constant460_outs),
    .data_valid (constant460_outs_valid),
    .data_ready (constant460_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br36_trueOut),
    .trueOut_valid (cond_br36_trueOut_valid),
    .trueOut_ready (cond_br36_trueOut_ready),
    .falseOut (cond_br36_falseOut),
    .falseOut_valid (cond_br36_falseOut_valid),
    .falseOut_ready (cond_br36_falseOut_ready)
  );

  sink #(.DATA_TYPE(15)) sink4(
    .ins (cond_br36_falseOut),
    .ins_valid (cond_br36_falseOut_valid),
    .ins_ready (cond_br36_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(15), .OUTPUT_TYPE(17)) extsi143(
    .ins (cond_br36_trueOut),
    .ins_valid (cond_br36_trueOut_valid),
    .ins_ready (cond_br36_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi143_outs),
    .outs_valid (extsi143_outs_valid),
    .outs_ready (extsi143_outs_ready)
  );

  cond_br #(.DATA_TYPE(12)) cond_br37(
    .condition (fork3_outs_2),
    .condition_valid (fork3_outs_2_valid),
    .condition_ready (fork3_outs_2_ready),
    .data (constant223_outs),
    .data_valid (constant223_outs_valid),
    .data_ready (constant223_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br37_trueOut),
    .trueOut_valid (cond_br37_trueOut_valid),
    .trueOut_ready (cond_br37_trueOut_ready),
    .falseOut (cond_br37_falseOut),
    .falseOut_valid (cond_br37_falseOut_valid),
    .falseOut_ready (cond_br37_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink5(
    .ins (cond_br37_falseOut),
    .ins_valid (cond_br37_falseOut_valid),
    .ins_ready (cond_br37_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br38(
    .condition (fork3_outs_0),
    .condition_valid (fork3_outs_0_valid),
    .condition_ready (fork3_outs_0_ready),
    .data (trunci13_outs),
    .data_valid (trunci13_outs_valid),
    .data_ready (trunci13_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br38_trueOut),
    .trueOut_valid (cond_br38_trueOut_valid),
    .trueOut_ready (cond_br38_trueOut_ready),
    .falseOut (cond_br38_falseOut),
    .falseOut_valid (cond_br38_falseOut_valid),
    .falseOut_ready (cond_br38_falseOut_ready)
  );

  cond_br_dataless cond_br39(
    .condition (fork3_outs_1),
    .condition_valid (fork3_outs_1_valid),
    .condition_ready (fork3_outs_1_ready),
    .data_valid (fork0_outs_7_valid),
    .data_ready (fork0_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br39_trueOut_valid),
    .trueOut_ready (cond_br39_trueOut_ready),
    .falseOut_valid (cond_br39_falseOut_valid),
    .falseOut_ready (cond_br39_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br40(
    .condition (fork3_outs_6),
    .condition_valid (fork3_outs_6_valid),
    .condition_ready (fork3_outs_6_ready),
    .data (fork2_outs_1),
    .data_valid (fork2_outs_1_valid),
    .data_ready (fork2_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br40_trueOut),
    .trueOut_valid (cond_br40_trueOut_valid),
    .trueOut_ready (cond_br40_trueOut_ready),
    .falseOut (cond_br40_falseOut),
    .falseOut_valid (cond_br40_falseOut_valid),
    .falseOut_ready (cond_br40_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink6(
    .ins (cond_br40_trueOut),
    .ins_valid (cond_br40_trueOut_valid),
    .ins_ready (cond_br40_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer2(
    .ins (cond_br40_falseOut),
    .ins_valid (cond_br40_falseOut_valid),
    .ins_ready (cond_br40_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer2_outs),
    .outs_valid (buffer2_outs_valid),
    .outs_ready (buffer2_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer3(
    .ins (buffer2_outs),
    .ins_valid (buffer2_outs_valid),
    .ins_ready (buffer2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer3_outs),
    .outs_valid (buffer3_outs_valid),
    .outs_ready (buffer3_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork4(
    .ins (buffer3_outs),
    .ins_valid (buffer3_outs_valid),
    .ins_ready (buffer3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork4_outs_1, fork4_outs_0}),
    .outs_valid ({fork4_outs_1_valid, fork4_outs_0_valid}),
    .outs_ready ({fork4_outs_1_ready, fork4_outs_0_ready})
  );

  oehb_dataless buffer4(
    .ins_valid (cond_br39_falseOut_valid),
    .ins_ready (cond_br39_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer4_outs_valid),
    .outs_ready (buffer4_outs_ready)
  );

  tehb_dataless buffer5(
    .ins_valid (buffer4_outs_valid),
    .ins_ready (buffer4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer5_outs_valid),
    .outs_ready (buffer5_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork5(
    .ins_valid (buffer5_outs_valid),
    .ins_ready (buffer5_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork5_outs_6_valid, fork5_outs_5_valid, fork5_outs_4_valid, fork5_outs_3_valid, fork5_outs_2_valid, fork5_outs_1_valid, fork5_outs_0_valid}),
    .outs_ready ({fork5_outs_6_ready, fork5_outs_5_ready, fork5_outs_4_ready, fork5_outs_3_ready, fork5_outs_2_ready, fork5_outs_1_ready, fork5_outs_0_ready})
  );

  handshake_constant_8 #(.DATA_WIDTH(34)) constant463(
    .ctrl_valid (fork5_outs_1_valid),
    .ctrl_ready (fork5_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant463_outs),
    .outs_valid (constant463_outs_valid),
    .outs_ready (constant463_outs_ready)
  );

  handshake_constant_9 #(.DATA_WIDTH(33)) constant231(
    .ctrl_valid (fork5_outs_5_valid),
    .ctrl_ready (fork5_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant231_outs),
    .outs_valid (constant231_outs_valid),
    .outs_ready (constant231_outs_ready)
  );

  handshake_constant_10 #(.DATA_WIDTH(27)) constant232(
    .ctrl_valid (fork5_outs_4_valid),
    .ctrl_ready (fork5_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant232_outs),
    .outs_valid (constant232_outs_valid),
    .outs_ready (constant232_outs_ready)
  );

  handshake_constant_11 #(.DATA_WIDTH(22)) constant233(
    .ctrl_valid (fork5_outs_3_valid),
    .ctrl_ready (fork5_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant233_outs),
    .outs_valid (constant233_outs_valid),
    .outs_ready (constant233_outs_ready)
  );

  handshake_constant_12 #(.DATA_WIDTH(16)) constant464(
    .ctrl_valid (fork5_outs_0_valid),
    .ctrl_ready (fork5_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant464_outs),
    .outs_valid (constant464_outs_valid),
    .outs_ready (constant464_outs_ready)
  );

  handshake_constant_13 #(.DATA_WIDTH(12)) constant235(
    .ctrl_valid (fork5_outs_2_valid),
    .ctrl_ready (fork5_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant235_outs),
    .outs_valid (constant235_outs_valid),
    .outs_ready (constant235_outs_ready)
  );

  source source2(
    .clk (clk),
    .rst (rst),
    .outs_valid (source2_outs_valid),
    .outs_ready (source2_outs_ready)
  );

  handshake_constant_14 #(.DATA_WIDTH(2)) constant465(
    .ctrl_valid (source2_outs_valid),
    .ctrl_ready (source2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant465_outs),
    .outs_valid (constant465_outs_valid),
    .outs_ready (constant465_outs_ready)
  );

  extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(5)) extsi144(
    .ins (constant465_outs),
    .ins_valid (constant465_outs_valid),
    .ins_ready (constant465_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi144_outs),
    .outs_valid (extsi144_outs_valid),
    .outs_ready (extsi144_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi1(
    .lhs (fork4_outs_0),
    .lhs_valid (fork4_outs_0_valid),
    .lhs_ready (fork4_outs_0_ready),
    .rhs (extsi144_outs),
    .rhs_valid (extsi144_outs_valid),
    .rhs_ready (extsi144_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi1_result),
    .result_valid (cmpi1_result_valid),
    .result_ready (cmpi1_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork6(
    .ins (cmpi1_result),
    .ins_valid (cmpi1_result_valid),
    .ins_ready (cmpi1_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork6_outs_8, fork6_outs_7, fork6_outs_6, fork6_outs_5, fork6_outs_4, fork6_outs_3, fork6_outs_2, fork6_outs_1, fork6_outs_0}),
    .outs_valid ({fork6_outs_8_valid, fork6_outs_7_valid, fork6_outs_6_valid, fork6_outs_5_valid, fork6_outs_4_valid, fork6_outs_3_valid, fork6_outs_2_valid, fork6_outs_1_valid, fork6_outs_0_valid}),
    .outs_ready ({fork6_outs_8_ready, fork6_outs_7_ready, fork6_outs_6_ready, fork6_outs_5_ready, fork6_outs_4_ready, fork6_outs_3_ready, fork6_outs_2_ready, fork6_outs_1_ready, fork6_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(34)) cond_br41(
    .condition (fork6_outs_7),
    .condition_valid (fork6_outs_7_valid),
    .condition_ready (fork6_outs_7_ready),
    .data (constant463_outs),
    .data_valid (constant463_outs_valid),
    .data_ready (constant463_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br41_trueOut),
    .trueOut_valid (cond_br41_trueOut_valid),
    .trueOut_ready (cond_br41_trueOut_ready),
    .falseOut (cond_br41_falseOut),
    .falseOut_valid (cond_br41_falseOut_valid),
    .falseOut_ready (cond_br41_falseOut_ready)
  );

  sink #(.DATA_TYPE(34)) sink8(
    .ins (cond_br41_falseOut),
    .ins_valid (cond_br41_falseOut_valid),
    .ins_ready (cond_br41_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(34), .OUTPUT_TYPE(37)) extsi145(
    .ins (cond_br41_trueOut),
    .ins_valid (cond_br41_trueOut_valid),
    .ins_ready (cond_br41_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi145_outs),
    .outs_valid (extsi145_outs_valid),
    .outs_ready (extsi145_outs_ready)
  );

  cond_br #(.DATA_TYPE(33)) cond_br42(
    .condition (fork6_outs_5),
    .condition_valid (fork6_outs_5_valid),
    .condition_ready (fork6_outs_5_ready),
    .data (constant231_outs),
    .data_valid (constant231_outs_valid),
    .data_ready (constant231_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br42_trueOut),
    .trueOut_valid (cond_br42_trueOut_valid),
    .trueOut_ready (cond_br42_trueOut_ready),
    .falseOut (cond_br42_falseOut),
    .falseOut_valid (cond_br42_falseOut_valid),
    .falseOut_ready (cond_br42_falseOut_ready)
  );

  sink #(.DATA_TYPE(33)) sink9(
    .ins (cond_br42_falseOut),
    .ins_valid (cond_br42_falseOut_valid),
    .ins_ready (cond_br42_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br43(
    .condition (fork6_outs_4),
    .condition_valid (fork6_outs_4_valid),
    .condition_ready (fork6_outs_4_ready),
    .data (constant232_outs),
    .data_valid (constant232_outs_valid),
    .data_ready (constant232_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br43_trueOut),
    .trueOut_valid (cond_br43_trueOut_valid),
    .trueOut_ready (cond_br43_trueOut_ready),
    .falseOut (cond_br43_falseOut),
    .falseOut_valid (cond_br43_falseOut_valid),
    .falseOut_ready (cond_br43_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink10(
    .ins (cond_br43_falseOut),
    .ins_valid (cond_br43_falseOut_valid),
    .ins_ready (cond_br43_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(22)) cond_br44(
    .condition (fork6_outs_3),
    .condition_valid (fork6_outs_3_valid),
    .condition_ready (fork6_outs_3_ready),
    .data (constant233_outs),
    .data_valid (constant233_outs_valid),
    .data_ready (constant233_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br44_trueOut),
    .trueOut_valid (cond_br44_trueOut_valid),
    .trueOut_ready (cond_br44_trueOut_ready),
    .falseOut (cond_br44_falseOut),
    .falseOut_valid (cond_br44_falseOut_valid),
    .falseOut_ready (cond_br44_falseOut_ready)
  );

  sink #(.DATA_TYPE(22)) sink11(
    .ins (cond_br44_falseOut),
    .ins_valid (cond_br44_falseOut_valid),
    .ins_ready (cond_br44_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(16)) cond_br45(
    .condition (fork6_outs_6),
    .condition_valid (fork6_outs_6_valid),
    .condition_ready (fork6_outs_6_ready),
    .data (constant464_outs),
    .data_valid (constant464_outs_valid),
    .data_ready (constant464_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br45_trueOut),
    .trueOut_valid (cond_br45_trueOut_valid),
    .trueOut_ready (cond_br45_trueOut_ready),
    .falseOut (cond_br45_falseOut),
    .falseOut_valid (cond_br45_falseOut_valid),
    .falseOut_ready (cond_br45_falseOut_ready)
  );

  sink #(.DATA_TYPE(16)) sink12(
    .ins (cond_br45_falseOut),
    .ins_valid (cond_br45_falseOut_valid),
    .ins_ready (cond_br45_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(16), .OUTPUT_TYPE(17)) extsi146(
    .ins (cond_br45_trueOut),
    .ins_valid (cond_br45_trueOut_valid),
    .ins_ready (cond_br45_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi146_outs),
    .outs_valid (extsi146_outs_valid),
    .outs_ready (extsi146_outs_ready)
  );

  cond_br #(.DATA_TYPE(12)) cond_br46(
    .condition (fork6_outs_2),
    .condition_valid (fork6_outs_2_valid),
    .condition_ready (fork6_outs_2_ready),
    .data (constant235_outs),
    .data_valid (constant235_outs_valid),
    .data_ready (constant235_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br46_trueOut),
    .trueOut_valid (cond_br46_trueOut_valid),
    .trueOut_ready (cond_br46_trueOut_ready),
    .falseOut (cond_br46_falseOut),
    .falseOut_valid (cond_br46_falseOut_valid),
    .falseOut_ready (cond_br46_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink13(
    .ins (cond_br46_falseOut),
    .ins_valid (cond_br46_falseOut_valid),
    .ins_ready (cond_br46_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer0(
    .ins (cond_br38_falseOut),
    .ins_valid (cond_br38_falseOut_valid),
    .ins_ready (cond_br38_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer0_outs),
    .outs_valid (buffer0_outs_valid),
    .outs_ready (buffer0_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer1(
    .ins (buffer0_outs),
    .ins_valid (buffer0_outs_valid),
    .ins_ready (buffer0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer1_outs),
    .outs_valid (buffer1_outs_valid),
    .outs_ready (buffer1_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br47(
    .condition (fork6_outs_0),
    .condition_valid (fork6_outs_0_valid),
    .condition_ready (fork6_outs_0_ready),
    .data (buffer1_outs),
    .data_valid (buffer1_outs_valid),
    .data_ready (buffer1_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br47_trueOut),
    .trueOut_valid (cond_br47_trueOut_valid),
    .trueOut_ready (cond_br47_trueOut_ready),
    .falseOut (cond_br47_falseOut),
    .falseOut_valid (cond_br47_falseOut_valid),
    .falseOut_ready (cond_br47_falseOut_ready)
  );

  cond_br_dataless cond_br48(
    .condition (fork6_outs_1),
    .condition_valid (fork6_outs_1_valid),
    .condition_ready (fork6_outs_1_ready),
    .data_valid (fork5_outs_6_valid),
    .data_ready (fork5_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br48_trueOut_valid),
    .trueOut_ready (cond_br48_trueOut_ready),
    .falseOut_valid (cond_br48_falseOut_valid),
    .falseOut_ready (cond_br48_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br49(
    .condition (fork6_outs_8),
    .condition_valid (fork6_outs_8_valid),
    .condition_ready (fork6_outs_8_ready),
    .data (fork4_outs_1),
    .data_valid (fork4_outs_1_valid),
    .data_ready (fork4_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br49_trueOut),
    .trueOut_valid (cond_br49_trueOut_valid),
    .trueOut_ready (cond_br49_trueOut_ready),
    .falseOut (cond_br49_falseOut),
    .falseOut_valid (cond_br49_falseOut_valid),
    .falseOut_ready (cond_br49_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink14(
    .ins (cond_br49_trueOut),
    .ins_valid (cond_br49_trueOut_valid),
    .ins_ready (cond_br49_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer8(
    .ins (cond_br49_falseOut),
    .ins_valid (cond_br49_falseOut_valid),
    .ins_ready (cond_br49_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer8_outs),
    .outs_valid (buffer8_outs_valid),
    .outs_ready (buffer8_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer9(
    .ins (buffer8_outs),
    .ins_valid (buffer8_outs_valid),
    .ins_ready (buffer8_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer9_outs),
    .outs_valid (buffer9_outs_valid),
    .outs_ready (buffer9_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork7(
    .ins (buffer9_outs),
    .ins_valid (buffer9_outs_valid),
    .ins_ready (buffer9_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork7_outs_1, fork7_outs_0}),
    .outs_valid ({fork7_outs_1_valid, fork7_outs_0_valid}),
    .outs_ready ({fork7_outs_1_ready, fork7_outs_0_ready})
  );

  oehb_dataless buffer10(
    .ins_valid (cond_br48_falseOut_valid),
    .ins_ready (cond_br48_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer10_outs_valid),
    .outs_ready (buffer10_outs_ready)
  );

  tehb_dataless buffer11(
    .ins_valid (buffer10_outs_valid),
    .ins_ready (buffer10_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer11_outs_valid),
    .outs_ready (buffer11_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork8(
    .ins_valid (buffer11_outs_valid),
    .ins_ready (buffer11_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork8_outs_6_valid, fork8_outs_5_valid, fork8_outs_4_valid, fork8_outs_3_valid, fork8_outs_2_valid, fork8_outs_1_valid, fork8_outs_0_valid}),
    .outs_ready ({fork8_outs_6_ready, fork8_outs_5_ready, fork8_outs_4_ready, fork8_outs_3_ready, fork8_outs_2_ready, fork8_outs_1_ready, fork8_outs_0_ready})
  );

  handshake_constant_15 #(.DATA_WIDTH(35)) constant466(
    .ctrl_valid (fork8_outs_0_valid),
    .ctrl_ready (fork8_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant466_outs),
    .outs_valid (constant466_outs_valid),
    .outs_ready (constant466_outs_ready)
  );

  handshake_constant_16 #(.DATA_WIDTH(33)) constant238(
    .ctrl_valid (fork8_outs_5_valid),
    .ctrl_ready (fork8_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant238_outs),
    .outs_valid (constant238_outs_valid),
    .outs_ready (constant238_outs_ready)
  );

  handshake_constant_17 #(.DATA_WIDTH(27)) constant239(
    .ctrl_valid (fork8_outs_4_valid),
    .ctrl_ready (fork8_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant239_outs),
    .outs_valid (constant239_outs_valid),
    .outs_ready (constant239_outs_ready)
  );

  handshake_constant_18 #(.DATA_WIDTH(22)) constant240(
    .ctrl_valid (fork8_outs_3_valid),
    .ctrl_ready (fork8_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant240_outs),
    .outs_valid (constant240_outs_valid),
    .outs_ready (constant240_outs_ready)
  );

  handshake_constant_19 #(.DATA_WIDTH(17)) constant241(
    .ctrl_valid (fork8_outs_2_valid),
    .ctrl_ready (fork8_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant241_outs),
    .outs_valid (constant241_outs_valid),
    .outs_ready (constant241_outs_ready)
  );

  handshake_constant_20 #(.DATA_WIDTH(12)) constant242(
    .ctrl_valid (fork8_outs_1_valid),
    .ctrl_ready (fork8_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant242_outs),
    .outs_valid (constant242_outs_valid),
    .outs_ready (constant242_outs_ready)
  );

  source source3(
    .clk (clk),
    .rst (rst),
    .outs_valid (source3_outs_valid),
    .outs_ready (source3_outs_ready)
  );

  handshake_constant_21 #(.DATA_WIDTH(3)) constant467(
    .ctrl_valid (source3_outs_valid),
    .ctrl_ready (source3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant467_outs),
    .outs_valid (constant467_outs_valid),
    .outs_ready (constant467_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(5)) extsi147(
    .ins (constant467_outs),
    .ins_valid (constant467_outs_valid),
    .ins_ready (constant467_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi147_outs),
    .outs_valid (extsi147_outs_valid),
    .outs_ready (extsi147_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi2(
    .lhs (fork7_outs_0),
    .lhs_valid (fork7_outs_0_valid),
    .lhs_ready (fork7_outs_0_ready),
    .rhs (extsi147_outs),
    .rhs_valid (extsi147_outs_valid),
    .rhs_ready (extsi147_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi2_result),
    .result_valid (cmpi2_result_valid),
    .result_ready (cmpi2_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork9(
    .ins (cmpi2_result),
    .ins_valid (cmpi2_result_valid),
    .ins_ready (cmpi2_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork9_outs_8, fork9_outs_7, fork9_outs_6, fork9_outs_5, fork9_outs_4, fork9_outs_3, fork9_outs_2, fork9_outs_1, fork9_outs_0}),
    .outs_valid ({fork9_outs_8_valid, fork9_outs_7_valid, fork9_outs_6_valid, fork9_outs_5_valid, fork9_outs_4_valid, fork9_outs_3_valid, fork9_outs_2_valid, fork9_outs_1_valid, fork9_outs_0_valid}),
    .outs_ready ({fork9_outs_8_ready, fork9_outs_7_ready, fork9_outs_6_ready, fork9_outs_5_ready, fork9_outs_4_ready, fork9_outs_3_ready, fork9_outs_2_ready, fork9_outs_1_ready, fork9_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(35)) cond_br50(
    .condition (fork9_outs_7),
    .condition_valid (fork9_outs_7_valid),
    .condition_ready (fork9_outs_7_ready),
    .data (constant466_outs),
    .data_valid (constant466_outs_valid),
    .data_ready (constant466_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br50_trueOut),
    .trueOut_valid (cond_br50_trueOut_valid),
    .trueOut_ready (cond_br50_trueOut_ready),
    .falseOut (cond_br50_falseOut),
    .falseOut_valid (cond_br50_falseOut_valid),
    .falseOut_ready (cond_br50_falseOut_ready)
  );

  sink #(.DATA_TYPE(35)) sink16(
    .ins (cond_br50_falseOut),
    .ins_valid (cond_br50_falseOut_valid),
    .ins_ready (cond_br50_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(35), .OUTPUT_TYPE(37)) extsi148(
    .ins (cond_br50_trueOut),
    .ins_valid (cond_br50_trueOut_valid),
    .ins_ready (cond_br50_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi148_outs),
    .outs_valid (extsi148_outs_valid),
    .outs_ready (extsi148_outs_ready)
  );

  cond_br #(.DATA_TYPE(33)) cond_br51(
    .condition (fork9_outs_6),
    .condition_valid (fork9_outs_6_valid),
    .condition_ready (fork9_outs_6_ready),
    .data (constant238_outs),
    .data_valid (constant238_outs_valid),
    .data_ready (constant238_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br51_trueOut),
    .trueOut_valid (cond_br51_trueOut_valid),
    .trueOut_ready (cond_br51_trueOut_ready),
    .falseOut (cond_br51_falseOut),
    .falseOut_valid (cond_br51_falseOut_valid),
    .falseOut_ready (cond_br51_falseOut_ready)
  );

  sink #(.DATA_TYPE(33)) sink17(
    .ins (cond_br51_falseOut),
    .ins_valid (cond_br51_falseOut_valid),
    .ins_ready (cond_br51_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br52(
    .condition (fork9_outs_5),
    .condition_valid (fork9_outs_5_valid),
    .condition_ready (fork9_outs_5_ready),
    .data (constant239_outs),
    .data_valid (constant239_outs_valid),
    .data_ready (constant239_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br52_trueOut),
    .trueOut_valid (cond_br52_trueOut_valid),
    .trueOut_ready (cond_br52_trueOut_ready),
    .falseOut (cond_br52_falseOut),
    .falseOut_valid (cond_br52_falseOut_valid),
    .falseOut_ready (cond_br52_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink18(
    .ins (cond_br52_falseOut),
    .ins_valid (cond_br52_falseOut_valid),
    .ins_ready (cond_br52_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(22)) cond_br53(
    .condition (fork9_outs_4),
    .condition_valid (fork9_outs_4_valid),
    .condition_ready (fork9_outs_4_ready),
    .data (constant240_outs),
    .data_valid (constant240_outs_valid),
    .data_ready (constant240_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br53_trueOut),
    .trueOut_valid (cond_br53_trueOut_valid),
    .trueOut_ready (cond_br53_trueOut_ready),
    .falseOut (cond_br53_falseOut),
    .falseOut_valid (cond_br53_falseOut_valid),
    .falseOut_ready (cond_br53_falseOut_ready)
  );

  sink #(.DATA_TYPE(22)) sink19(
    .ins (cond_br53_falseOut),
    .ins_valid (cond_br53_falseOut_valid),
    .ins_ready (cond_br53_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(17)) cond_br54(
    .condition (fork9_outs_3),
    .condition_valid (fork9_outs_3_valid),
    .condition_ready (fork9_outs_3_ready),
    .data (constant241_outs),
    .data_valid (constant241_outs_valid),
    .data_ready (constant241_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br54_trueOut),
    .trueOut_valid (cond_br54_trueOut_valid),
    .trueOut_ready (cond_br54_trueOut_ready),
    .falseOut (cond_br54_falseOut),
    .falseOut_valid (cond_br54_falseOut_valid),
    .falseOut_ready (cond_br54_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink20(
    .ins (cond_br54_falseOut),
    .ins_valid (cond_br54_falseOut_valid),
    .ins_ready (cond_br54_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br55(
    .condition (fork9_outs_2),
    .condition_valid (fork9_outs_2_valid),
    .condition_ready (fork9_outs_2_ready),
    .data (constant242_outs),
    .data_valid (constant242_outs_valid),
    .data_ready (constant242_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br55_trueOut),
    .trueOut_valid (cond_br55_trueOut_valid),
    .trueOut_ready (cond_br55_trueOut_ready),
    .falseOut (cond_br55_falseOut),
    .falseOut_valid (cond_br55_falseOut_valid),
    .falseOut_ready (cond_br55_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink21(
    .ins (cond_br55_falseOut),
    .ins_valid (cond_br55_falseOut_valid),
    .ins_ready (cond_br55_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer6(
    .ins (cond_br47_falseOut),
    .ins_valid (cond_br47_falseOut_valid),
    .ins_ready (cond_br47_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer6_outs),
    .outs_valid (buffer6_outs_valid),
    .outs_ready (buffer6_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer7(
    .ins (buffer6_outs),
    .ins_valid (buffer6_outs_valid),
    .ins_ready (buffer6_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer7_outs),
    .outs_valid (buffer7_outs_valid),
    .outs_ready (buffer7_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br56(
    .condition (fork9_outs_0),
    .condition_valid (fork9_outs_0_valid),
    .condition_ready (fork9_outs_0_ready),
    .data (buffer7_outs),
    .data_valid (buffer7_outs_valid),
    .data_ready (buffer7_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br56_trueOut),
    .trueOut_valid (cond_br56_trueOut_valid),
    .trueOut_ready (cond_br56_trueOut_ready),
    .falseOut (cond_br56_falseOut),
    .falseOut_valid (cond_br56_falseOut_valid),
    .falseOut_ready (cond_br56_falseOut_ready)
  );

  cond_br_dataless cond_br57(
    .condition (fork9_outs_1),
    .condition_valid (fork9_outs_1_valid),
    .condition_ready (fork9_outs_1_ready),
    .data_valid (fork8_outs_6_valid),
    .data_ready (fork8_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br57_trueOut_valid),
    .trueOut_ready (cond_br57_trueOut_ready),
    .falseOut_valid (cond_br57_falseOut_valid),
    .falseOut_ready (cond_br57_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br58(
    .condition (fork9_outs_8),
    .condition_valid (fork9_outs_8_valid),
    .condition_ready (fork9_outs_8_ready),
    .data (fork7_outs_1),
    .data_valid (fork7_outs_1_valid),
    .data_ready (fork7_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br58_trueOut),
    .trueOut_valid (cond_br58_trueOut_valid),
    .trueOut_ready (cond_br58_trueOut_ready),
    .falseOut (cond_br58_falseOut),
    .falseOut_valid (cond_br58_falseOut_valid),
    .falseOut_ready (cond_br58_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink22(
    .ins (cond_br58_trueOut),
    .ins_valid (cond_br58_trueOut_valid),
    .ins_ready (cond_br58_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer14(
    .ins (cond_br58_falseOut),
    .ins_valid (cond_br58_falseOut_valid),
    .ins_ready (cond_br58_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer14_outs),
    .outs_valid (buffer14_outs_valid),
    .outs_ready (buffer14_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer15(
    .ins (buffer14_outs),
    .ins_valid (buffer14_outs_valid),
    .ins_ready (buffer14_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer15_outs),
    .outs_valid (buffer15_outs_valid),
    .outs_ready (buffer15_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork10(
    .ins (buffer15_outs),
    .ins_valid (buffer15_outs_valid),
    .ins_ready (buffer15_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork10_outs_1, fork10_outs_0}),
    .outs_valid ({fork10_outs_1_valid, fork10_outs_0_valid}),
    .outs_ready ({fork10_outs_1_ready, fork10_outs_0_ready})
  );

  oehb_dataless buffer16(
    .ins_valid (cond_br57_falseOut_valid),
    .ins_ready (cond_br57_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer16_outs_valid),
    .outs_ready (buffer16_outs_ready)
  );

  tehb_dataless buffer17(
    .ins_valid (buffer16_outs_valid),
    .ins_ready (buffer16_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer17_outs_valid),
    .outs_ready (buffer17_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork11(
    .ins_valid (buffer17_outs_valid),
    .ins_ready (buffer17_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork11_outs_6_valid, fork11_outs_5_valid, fork11_outs_4_valid, fork11_outs_3_valid, fork11_outs_2_valid, fork11_outs_1_valid, fork11_outs_0_valid}),
    .outs_ready ({fork11_outs_6_ready, fork11_outs_5_ready, fork11_outs_4_ready, fork11_outs_3_ready, fork11_outs_2_ready, fork11_outs_1_ready, fork11_outs_0_ready})
  );

  handshake_constant_22 #(.DATA_WIDTH(36)) constant468(
    .ctrl_valid (fork11_outs_1_valid),
    .ctrl_ready (fork11_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant468_outs),
    .outs_valid (constant468_outs_valid),
    .outs_ready (constant468_outs_ready)
  );

  handshake_constant_23 #(.DATA_WIDTH(33)) constant245(
    .ctrl_valid (fork11_outs_5_valid),
    .ctrl_ready (fork11_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant245_outs),
    .outs_valid (constant245_outs_valid),
    .outs_ready (constant245_outs_ready)
  );

  handshake_constant_24 #(.DATA_WIDTH(27)) constant246(
    .ctrl_valid (fork11_outs_4_valid),
    .ctrl_ready (fork11_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant246_outs),
    .outs_valid (constant246_outs_valid),
    .outs_ready (constant246_outs_ready)
  );

  handshake_constant_25 #(.DATA_WIDTH(22)) constant247(
    .ctrl_valid (fork11_outs_3_valid),
    .ctrl_ready (fork11_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant247_outs),
    .outs_valid (constant247_outs_valid),
    .outs_ready (constant247_outs_ready)
  );

  handshake_constant_26 #(.DATA_WIDTH(17)) constant248(
    .ctrl_valid (fork11_outs_2_valid),
    .ctrl_ready (fork11_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant248_outs),
    .outs_valid (constant248_outs_valid),
    .outs_ready (constant248_outs_ready)
  );

  handshake_constant_27 #(.DATA_WIDTH(11)) constant469(
    .ctrl_valid (fork11_outs_0_valid),
    .ctrl_ready (fork11_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant469_outs),
    .outs_valid (constant469_outs_valid),
    .outs_ready (constant469_outs_ready)
  );

  source source4(
    .clk (clk),
    .rst (rst),
    .outs_valid (source4_outs_valid),
    .outs_ready (source4_outs_ready)
  );

  handshake_constant_28 #(.DATA_WIDTH(3)) constant470(
    .ctrl_valid (source4_outs_valid),
    .ctrl_ready (source4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant470_outs),
    .outs_valid (constant470_outs_valid),
    .outs_ready (constant470_outs_ready)
  );

  extsi #(.INPUT_TYPE(3), .OUTPUT_TYPE(5)) extsi149(
    .ins (constant470_outs),
    .ins_valid (constant470_outs_valid),
    .ins_ready (constant470_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi149_outs),
    .outs_valid (extsi149_outs_valid),
    .outs_ready (extsi149_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi3(
    .lhs (fork10_outs_0),
    .lhs_valid (fork10_outs_0_valid),
    .lhs_ready (fork10_outs_0_ready),
    .rhs (extsi149_outs),
    .rhs_valid (extsi149_outs_valid),
    .rhs_ready (extsi149_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi3_result),
    .result_valid (cmpi3_result_valid),
    .result_ready (cmpi3_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork12(
    .ins (cmpi3_result),
    .ins_valid (cmpi3_result_valid),
    .ins_ready (cmpi3_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork12_outs_8, fork12_outs_7, fork12_outs_6, fork12_outs_5, fork12_outs_4, fork12_outs_3, fork12_outs_2, fork12_outs_1, fork12_outs_0}),
    .outs_valid ({fork12_outs_8_valid, fork12_outs_7_valid, fork12_outs_6_valid, fork12_outs_5_valid, fork12_outs_4_valid, fork12_outs_3_valid, fork12_outs_2_valid, fork12_outs_1_valid, fork12_outs_0_valid}),
    .outs_ready ({fork12_outs_8_ready, fork12_outs_7_ready, fork12_outs_6_ready, fork12_outs_5_ready, fork12_outs_4_ready, fork12_outs_3_ready, fork12_outs_2_ready, fork12_outs_1_ready, fork12_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(36)) cond_br59(
    .condition (fork12_outs_7),
    .condition_valid (fork12_outs_7_valid),
    .condition_ready (fork12_outs_7_ready),
    .data (constant468_outs),
    .data_valid (constant468_outs_valid),
    .data_ready (constant468_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br59_trueOut),
    .trueOut_valid (cond_br59_trueOut_valid),
    .trueOut_ready (cond_br59_trueOut_ready),
    .falseOut (cond_br59_falseOut),
    .falseOut_valid (cond_br59_falseOut_valid),
    .falseOut_ready (cond_br59_falseOut_ready)
  );

  sink #(.DATA_TYPE(36)) sink24(
    .ins (cond_br59_falseOut),
    .ins_valid (cond_br59_falseOut_valid),
    .ins_ready (cond_br59_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(36), .OUTPUT_TYPE(37)) extsi150(
    .ins (cond_br59_trueOut),
    .ins_valid (cond_br59_trueOut_valid),
    .ins_ready (cond_br59_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi150_outs),
    .outs_valid (extsi150_outs_valid),
    .outs_ready (extsi150_outs_ready)
  );

  cond_br #(.DATA_TYPE(33)) cond_br60(
    .condition (fork12_outs_5),
    .condition_valid (fork12_outs_5_valid),
    .condition_ready (fork12_outs_5_ready),
    .data (constant245_outs),
    .data_valid (constant245_outs_valid),
    .data_ready (constant245_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br60_trueOut),
    .trueOut_valid (cond_br60_trueOut_valid),
    .trueOut_ready (cond_br60_trueOut_ready),
    .falseOut (cond_br60_falseOut),
    .falseOut_valid (cond_br60_falseOut_valid),
    .falseOut_ready (cond_br60_falseOut_ready)
  );

  sink #(.DATA_TYPE(33)) sink25(
    .ins (cond_br60_falseOut),
    .ins_valid (cond_br60_falseOut_valid),
    .ins_ready (cond_br60_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br61(
    .condition (fork12_outs_4),
    .condition_valid (fork12_outs_4_valid),
    .condition_ready (fork12_outs_4_ready),
    .data (constant246_outs),
    .data_valid (constant246_outs_valid),
    .data_ready (constant246_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br61_trueOut),
    .trueOut_valid (cond_br61_trueOut_valid),
    .trueOut_ready (cond_br61_trueOut_ready),
    .falseOut (cond_br61_falseOut),
    .falseOut_valid (cond_br61_falseOut_valid),
    .falseOut_ready (cond_br61_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink26(
    .ins (cond_br61_falseOut),
    .ins_valid (cond_br61_falseOut_valid),
    .ins_ready (cond_br61_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(22)) cond_br62(
    .condition (fork12_outs_3),
    .condition_valid (fork12_outs_3_valid),
    .condition_ready (fork12_outs_3_ready),
    .data (constant247_outs),
    .data_valid (constant247_outs_valid),
    .data_ready (constant247_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br62_trueOut),
    .trueOut_valid (cond_br62_trueOut_valid),
    .trueOut_ready (cond_br62_trueOut_ready),
    .falseOut (cond_br62_falseOut),
    .falseOut_valid (cond_br62_falseOut_valid),
    .falseOut_ready (cond_br62_falseOut_ready)
  );

  sink #(.DATA_TYPE(22)) sink27(
    .ins (cond_br62_falseOut),
    .ins_valid (cond_br62_falseOut_valid),
    .ins_ready (cond_br62_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(17)) cond_br63(
    .condition (fork12_outs_2),
    .condition_valid (fork12_outs_2_valid),
    .condition_ready (fork12_outs_2_ready),
    .data (constant248_outs),
    .data_valid (constant248_outs_valid),
    .data_ready (constant248_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br63_trueOut),
    .trueOut_valid (cond_br63_trueOut_valid),
    .trueOut_ready (cond_br63_trueOut_ready),
    .falseOut (cond_br63_falseOut),
    .falseOut_valid (cond_br63_falseOut_valid),
    .falseOut_ready (cond_br63_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink28(
    .ins (cond_br63_falseOut),
    .ins_valid (cond_br63_falseOut_valid),
    .ins_ready (cond_br63_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(11)) cond_br64(
    .condition (fork12_outs_6),
    .condition_valid (fork12_outs_6_valid),
    .condition_ready (fork12_outs_6_ready),
    .data (constant469_outs),
    .data_valid (constant469_outs_valid),
    .data_ready (constant469_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br64_trueOut),
    .trueOut_valid (cond_br64_trueOut_valid),
    .trueOut_ready (cond_br64_trueOut_ready),
    .falseOut (cond_br64_falseOut),
    .falseOut_valid (cond_br64_falseOut_valid),
    .falseOut_ready (cond_br64_falseOut_ready)
  );

  sink #(.DATA_TYPE(11)) sink29(
    .ins (cond_br64_falseOut),
    .ins_valid (cond_br64_falseOut_valid),
    .ins_ready (cond_br64_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(11), .OUTPUT_TYPE(12)) extsi151(
    .ins (cond_br64_trueOut),
    .ins_valid (cond_br64_trueOut_valid),
    .ins_ready (cond_br64_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi151_outs),
    .outs_valid (extsi151_outs_valid),
    .outs_ready (extsi151_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer12(
    .ins (cond_br56_falseOut),
    .ins_valid (cond_br56_falseOut_valid),
    .ins_ready (cond_br56_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer12_outs),
    .outs_valid (buffer12_outs_valid),
    .outs_ready (buffer12_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer13(
    .ins (buffer12_outs),
    .ins_valid (buffer12_outs_valid),
    .ins_ready (buffer12_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer13_outs),
    .outs_valid (buffer13_outs_valid),
    .outs_ready (buffer13_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br65(
    .condition (fork12_outs_0),
    .condition_valid (fork12_outs_0_valid),
    .condition_ready (fork12_outs_0_ready),
    .data (buffer13_outs),
    .data_valid (buffer13_outs_valid),
    .data_ready (buffer13_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br65_trueOut),
    .trueOut_valid (cond_br65_trueOut_valid),
    .trueOut_ready (cond_br65_trueOut_ready),
    .falseOut (cond_br65_falseOut),
    .falseOut_valid (cond_br65_falseOut_valid),
    .falseOut_ready (cond_br65_falseOut_ready)
  );

  cond_br_dataless cond_br66(
    .condition (fork12_outs_1),
    .condition_valid (fork12_outs_1_valid),
    .condition_ready (fork12_outs_1_ready),
    .data_valid (fork11_outs_6_valid),
    .data_ready (fork11_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br66_trueOut_valid),
    .trueOut_ready (cond_br66_trueOut_ready),
    .falseOut_valid (cond_br66_falseOut_valid),
    .falseOut_ready (cond_br66_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br67(
    .condition (fork12_outs_8),
    .condition_valid (fork12_outs_8_valid),
    .condition_ready (fork12_outs_8_ready),
    .data (fork10_outs_1),
    .data_valid (fork10_outs_1_valid),
    .data_ready (fork10_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br67_trueOut),
    .trueOut_valid (cond_br67_trueOut_valid),
    .trueOut_ready (cond_br67_trueOut_ready),
    .falseOut (cond_br67_falseOut),
    .falseOut_valid (cond_br67_falseOut_valid),
    .falseOut_ready (cond_br67_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink30(
    .ins (cond_br67_trueOut),
    .ins_valid (cond_br67_trueOut_valid),
    .ins_ready (cond_br67_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer20(
    .ins (cond_br67_falseOut),
    .ins_valid (cond_br67_falseOut_valid),
    .ins_ready (cond_br67_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer20_outs),
    .outs_valid (buffer20_outs_valid),
    .outs_ready (buffer20_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer21(
    .ins (buffer20_outs),
    .ins_valid (buffer20_outs_valid),
    .ins_ready (buffer20_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer21_outs),
    .outs_valid (buffer21_outs_valid),
    .outs_ready (buffer21_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork13(
    .ins (buffer21_outs),
    .ins_valid (buffer21_outs_valid),
    .ins_ready (buffer21_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork13_outs_1, fork13_outs_0}),
    .outs_valid ({fork13_outs_1_valid, fork13_outs_0_valid}),
    .outs_ready ({fork13_outs_1_ready, fork13_outs_0_ready})
  );

  oehb_dataless buffer22(
    .ins_valid (cond_br66_falseOut_valid),
    .ins_ready (cond_br66_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer22_outs_valid),
    .outs_ready (buffer22_outs_ready)
  );

  tehb_dataless buffer23(
    .ins_valid (buffer22_outs_valid),
    .ins_ready (buffer22_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer23_outs_valid),
    .outs_ready (buffer23_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork14(
    .ins_valid (buffer23_outs_valid),
    .ins_ready (buffer23_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork14_outs_6_valid, fork14_outs_5_valid, fork14_outs_4_valid, fork14_outs_3_valid, fork14_outs_2_valid, fork14_outs_1_valid, fork14_outs_0_valid}),
    .outs_ready ({fork14_outs_6_ready, fork14_outs_5_ready, fork14_outs_4_ready, fork14_outs_3_ready, fork14_outs_2_ready, fork14_outs_1_ready, fork14_outs_0_ready})
  );

  handshake_constant_29 #(.DATA_WIDTH(36)) constant471(
    .ctrl_valid (fork14_outs_0_valid),
    .ctrl_ready (fork14_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant471_outs),
    .outs_valid (constant471_outs_valid),
    .outs_ready (constant471_outs_ready)
  );

  handshake_constant_30 #(.DATA_WIDTH(33)) constant252(
    .ctrl_valid (fork14_outs_5_valid),
    .ctrl_ready (fork14_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant252_outs),
    .outs_valid (constant252_outs_valid),
    .outs_ready (constant252_outs_ready)
  );

  handshake_constant_31 #(.DATA_WIDTH(27)) constant253(
    .ctrl_valid (fork14_outs_4_valid),
    .ctrl_ready (fork14_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant253_outs),
    .outs_valid (constant253_outs_valid),
    .outs_ready (constant253_outs_ready)
  );

  handshake_constant_32 #(.DATA_WIDTH(22)) constant254(
    .ctrl_valid (fork14_outs_3_valid),
    .ctrl_ready (fork14_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant254_outs),
    .outs_valid (constant254_outs_valid),
    .outs_ready (constant254_outs_ready)
  );

  handshake_constant_33 #(.DATA_WIDTH(17)) constant255(
    .ctrl_valid (fork14_outs_2_valid),
    .ctrl_ready (fork14_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant255_outs),
    .outs_valid (constant255_outs_valid),
    .outs_ready (constant255_outs_ready)
  );

  handshake_constant_34 #(.DATA_WIDTH(12)) constant256(
    .ctrl_valid (fork14_outs_1_valid),
    .ctrl_ready (fork14_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant256_outs),
    .outs_valid (constant256_outs_valid),
    .outs_ready (constant256_outs_ready)
  );

  source source5(
    .clk (clk),
    .rst (rst),
    .outs_valid (source5_outs_valid),
    .outs_ready (source5_outs_ready)
  );

  handshake_constant_35 #(.DATA_WIDTH(4)) constant472(
    .ctrl_valid (source5_outs_valid),
    .ctrl_ready (source5_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant472_outs),
    .outs_valid (constant472_outs_valid),
    .outs_ready (constant472_outs_ready)
  );

  extsi #(.INPUT_TYPE(4), .OUTPUT_TYPE(5)) extsi152(
    .ins (constant472_outs),
    .ins_valid (constant472_outs_valid),
    .ins_ready (constant472_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi152_outs),
    .outs_valid (extsi152_outs_valid),
    .outs_ready (extsi152_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi4(
    .lhs (fork13_outs_0),
    .lhs_valid (fork13_outs_0_valid),
    .lhs_ready (fork13_outs_0_ready),
    .rhs (extsi152_outs),
    .rhs_valid (extsi152_outs_valid),
    .rhs_ready (extsi152_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi4_result),
    .result_valid (cmpi4_result_valid),
    .result_ready (cmpi4_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork15(
    .ins (cmpi4_result),
    .ins_valid (cmpi4_result_valid),
    .ins_ready (cmpi4_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork15_outs_8, fork15_outs_7, fork15_outs_6, fork15_outs_5, fork15_outs_4, fork15_outs_3, fork15_outs_2, fork15_outs_1, fork15_outs_0}),
    .outs_valid ({fork15_outs_8_valid, fork15_outs_7_valid, fork15_outs_6_valid, fork15_outs_5_valid, fork15_outs_4_valid, fork15_outs_3_valid, fork15_outs_2_valid, fork15_outs_1_valid, fork15_outs_0_valid}),
    .outs_ready ({fork15_outs_8_ready, fork15_outs_7_ready, fork15_outs_6_ready, fork15_outs_5_ready, fork15_outs_4_ready, fork15_outs_3_ready, fork15_outs_2_ready, fork15_outs_1_ready, fork15_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(36)) cond_br68(
    .condition (fork15_outs_7),
    .condition_valid (fork15_outs_7_valid),
    .condition_ready (fork15_outs_7_ready),
    .data (constant471_outs),
    .data_valid (constant471_outs_valid),
    .data_ready (constant471_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br68_trueOut),
    .trueOut_valid (cond_br68_trueOut_valid),
    .trueOut_ready (cond_br68_trueOut_ready),
    .falseOut (cond_br68_falseOut),
    .falseOut_valid (cond_br68_falseOut_valid),
    .falseOut_ready (cond_br68_falseOut_ready)
  );

  sink #(.DATA_TYPE(36)) sink32(
    .ins (cond_br68_falseOut),
    .ins_valid (cond_br68_falseOut_valid),
    .ins_ready (cond_br68_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(36), .OUTPUT_TYPE(37)) extsi153(
    .ins (cond_br68_trueOut),
    .ins_valid (cond_br68_trueOut_valid),
    .ins_ready (cond_br68_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi153_outs),
    .outs_valid (extsi153_outs_valid),
    .outs_ready (extsi153_outs_ready)
  );

  cond_br #(.DATA_TYPE(33)) cond_br69(
    .condition (fork15_outs_6),
    .condition_valid (fork15_outs_6_valid),
    .condition_ready (fork15_outs_6_ready),
    .data (constant252_outs),
    .data_valid (constant252_outs_valid),
    .data_ready (constant252_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br69_trueOut),
    .trueOut_valid (cond_br69_trueOut_valid),
    .trueOut_ready (cond_br69_trueOut_ready),
    .falseOut (cond_br69_falseOut),
    .falseOut_valid (cond_br69_falseOut_valid),
    .falseOut_ready (cond_br69_falseOut_ready)
  );

  sink #(.DATA_TYPE(33)) sink33(
    .ins (cond_br69_falseOut),
    .ins_valid (cond_br69_falseOut_valid),
    .ins_ready (cond_br69_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br70(
    .condition (fork15_outs_5),
    .condition_valid (fork15_outs_5_valid),
    .condition_ready (fork15_outs_5_ready),
    .data (constant253_outs),
    .data_valid (constant253_outs_valid),
    .data_ready (constant253_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br70_trueOut),
    .trueOut_valid (cond_br70_trueOut_valid),
    .trueOut_ready (cond_br70_trueOut_ready),
    .falseOut (cond_br70_falseOut),
    .falseOut_valid (cond_br70_falseOut_valid),
    .falseOut_ready (cond_br70_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink34(
    .ins (cond_br70_falseOut),
    .ins_valid (cond_br70_falseOut_valid),
    .ins_ready (cond_br70_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(22)) cond_br71(
    .condition (fork15_outs_4),
    .condition_valid (fork15_outs_4_valid),
    .condition_ready (fork15_outs_4_ready),
    .data (constant254_outs),
    .data_valid (constant254_outs_valid),
    .data_ready (constant254_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br71_trueOut),
    .trueOut_valid (cond_br71_trueOut_valid),
    .trueOut_ready (cond_br71_trueOut_ready),
    .falseOut (cond_br71_falseOut),
    .falseOut_valid (cond_br71_falseOut_valid),
    .falseOut_ready (cond_br71_falseOut_ready)
  );

  sink #(.DATA_TYPE(22)) sink35(
    .ins (cond_br71_falseOut),
    .ins_valid (cond_br71_falseOut_valid),
    .ins_ready (cond_br71_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(17)) cond_br72(
    .condition (fork15_outs_3),
    .condition_valid (fork15_outs_3_valid),
    .condition_ready (fork15_outs_3_ready),
    .data (constant255_outs),
    .data_valid (constant255_outs_valid),
    .data_ready (constant255_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br72_trueOut),
    .trueOut_valid (cond_br72_trueOut_valid),
    .trueOut_ready (cond_br72_trueOut_ready),
    .falseOut (cond_br72_falseOut),
    .falseOut_valid (cond_br72_falseOut_valid),
    .falseOut_ready (cond_br72_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink36(
    .ins (cond_br72_falseOut),
    .ins_valid (cond_br72_falseOut_valid),
    .ins_ready (cond_br72_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br73(
    .condition (fork15_outs_2),
    .condition_valid (fork15_outs_2_valid),
    .condition_ready (fork15_outs_2_ready),
    .data (constant256_outs),
    .data_valid (constant256_outs_valid),
    .data_ready (constant256_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br73_trueOut),
    .trueOut_valid (cond_br73_trueOut_valid),
    .trueOut_ready (cond_br73_trueOut_ready),
    .falseOut (cond_br73_falseOut),
    .falseOut_valid (cond_br73_falseOut_valid),
    .falseOut_ready (cond_br73_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink37(
    .ins (cond_br73_falseOut),
    .ins_valid (cond_br73_falseOut_valid),
    .ins_ready (cond_br73_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer18(
    .ins (cond_br65_falseOut),
    .ins_valid (cond_br65_falseOut_valid),
    .ins_ready (cond_br65_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer18_outs),
    .outs_valid (buffer18_outs_valid),
    .outs_ready (buffer18_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer19(
    .ins (buffer18_outs),
    .ins_valid (buffer18_outs_valid),
    .ins_ready (buffer18_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer19_outs),
    .outs_valid (buffer19_outs_valid),
    .outs_ready (buffer19_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br74(
    .condition (fork15_outs_0),
    .condition_valid (fork15_outs_0_valid),
    .condition_ready (fork15_outs_0_ready),
    .data (buffer19_outs),
    .data_valid (buffer19_outs_valid),
    .data_ready (buffer19_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br74_trueOut),
    .trueOut_valid (cond_br74_trueOut_valid),
    .trueOut_ready (cond_br74_trueOut_ready),
    .falseOut (cond_br74_falseOut),
    .falseOut_valid (cond_br74_falseOut_valid),
    .falseOut_ready (cond_br74_falseOut_ready)
  );

  cond_br_dataless cond_br75(
    .condition (fork15_outs_1),
    .condition_valid (fork15_outs_1_valid),
    .condition_ready (fork15_outs_1_ready),
    .data_valid (fork14_outs_6_valid),
    .data_ready (fork14_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br75_trueOut_valid),
    .trueOut_ready (cond_br75_trueOut_ready),
    .falseOut_valid (cond_br75_falseOut_valid),
    .falseOut_ready (cond_br75_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br76(
    .condition (fork15_outs_8),
    .condition_valid (fork15_outs_8_valid),
    .condition_ready (fork15_outs_8_ready),
    .data (fork13_outs_1),
    .data_valid (fork13_outs_1_valid),
    .data_ready (fork13_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br76_trueOut),
    .trueOut_valid (cond_br76_trueOut_valid),
    .trueOut_ready (cond_br76_trueOut_ready),
    .falseOut (cond_br76_falseOut),
    .falseOut_valid (cond_br76_falseOut_valid),
    .falseOut_ready (cond_br76_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink38(
    .ins (cond_br76_trueOut),
    .ins_valid (cond_br76_trueOut_valid),
    .ins_ready (cond_br76_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer26(
    .ins (cond_br76_falseOut),
    .ins_valid (cond_br76_falseOut_valid),
    .ins_ready (cond_br76_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer26_outs),
    .outs_valid (buffer26_outs_valid),
    .outs_ready (buffer26_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer27(
    .ins (buffer26_outs),
    .ins_valid (buffer26_outs_valid),
    .ins_ready (buffer26_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer27_outs),
    .outs_valid (buffer27_outs_valid),
    .outs_ready (buffer27_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork16(
    .ins (buffer27_outs),
    .ins_valid (buffer27_outs_valid),
    .ins_ready (buffer27_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork16_outs_1, fork16_outs_0}),
    .outs_valid ({fork16_outs_1_valid, fork16_outs_0_valid}),
    .outs_ready ({fork16_outs_1_ready, fork16_outs_0_ready})
  );

  oehb_dataless buffer28(
    .ins_valid (cond_br75_falseOut_valid),
    .ins_ready (cond_br75_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer28_outs_valid),
    .outs_ready (buffer28_outs_ready)
  );

  tehb_dataless buffer29(
    .ins_valid (buffer28_outs_valid),
    .ins_ready (buffer28_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer29_outs_valid),
    .outs_ready (buffer29_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork17(
    .ins_valid (buffer29_outs_valid),
    .ins_ready (buffer29_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork17_outs_6_valid, fork17_outs_5_valid, fork17_outs_4_valid, fork17_outs_3_valid, fork17_outs_2_valid, fork17_outs_1_valid, fork17_outs_0_valid}),
    .outs_ready ({fork17_outs_6_ready, fork17_outs_5_ready, fork17_outs_4_ready, fork17_outs_3_ready, fork17_outs_2_ready, fork17_outs_1_ready, fork17_outs_0_ready})
  );

  handshake_constant_36 #(.DATA_WIDTH(36)) constant473(
    .ctrl_valid (fork17_outs_0_valid),
    .ctrl_ready (fork17_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant473_outs),
    .outs_valid (constant473_outs_valid),
    .outs_ready (constant473_outs_ready)
  );

  handshake_constant_37 #(.DATA_WIDTH(33)) constant259(
    .ctrl_valid (fork17_outs_5_valid),
    .ctrl_ready (fork17_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant259_outs),
    .outs_valid (constant259_outs_valid),
    .outs_ready (constant259_outs_ready)
  );

  handshake_constant_38 #(.DATA_WIDTH(27)) constant260(
    .ctrl_valid (fork17_outs_4_valid),
    .ctrl_ready (fork17_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant260_outs),
    .outs_valid (constant260_outs_valid),
    .outs_ready (constant260_outs_ready)
  );

  handshake_constant_39 #(.DATA_WIDTH(22)) constant261(
    .ctrl_valid (fork17_outs_3_valid),
    .ctrl_ready (fork17_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant261_outs),
    .outs_valid (constant261_outs_valid),
    .outs_ready (constant261_outs_ready)
  );

  handshake_constant_40 #(.DATA_WIDTH(17)) constant262(
    .ctrl_valid (fork17_outs_2_valid),
    .ctrl_ready (fork17_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant262_outs),
    .outs_valid (constant262_outs_valid),
    .outs_ready (constant262_outs_ready)
  );

  handshake_constant_41 #(.DATA_WIDTH(12)) constant263(
    .ctrl_valid (fork17_outs_1_valid),
    .ctrl_ready (fork17_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant263_outs),
    .outs_valid (constant263_outs_valid),
    .outs_ready (constant263_outs_ready)
  );

  source source6(
    .clk (clk),
    .rst (rst),
    .outs_valid (source6_outs_valid),
    .outs_ready (source6_outs_ready)
  );

  handshake_constant_42 #(.DATA_WIDTH(4)) constant474(
    .ctrl_valid (source6_outs_valid),
    .ctrl_ready (source6_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant474_outs),
    .outs_valid (constant474_outs_valid),
    .outs_ready (constant474_outs_ready)
  );

  extsi #(.INPUT_TYPE(4), .OUTPUT_TYPE(5)) extsi154(
    .ins (constant474_outs),
    .ins_valid (constant474_outs_valid),
    .ins_ready (constant474_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi154_outs),
    .outs_valid (extsi154_outs_valid),
    .outs_ready (extsi154_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi5(
    .lhs (fork16_outs_0),
    .lhs_valid (fork16_outs_0_valid),
    .lhs_ready (fork16_outs_0_ready),
    .rhs (extsi154_outs),
    .rhs_valid (extsi154_outs_valid),
    .rhs_ready (extsi154_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi5_result),
    .result_valid (cmpi5_result_valid),
    .result_ready (cmpi5_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork18(
    .ins (cmpi5_result),
    .ins_valid (cmpi5_result_valid),
    .ins_ready (cmpi5_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork18_outs_8, fork18_outs_7, fork18_outs_6, fork18_outs_5, fork18_outs_4, fork18_outs_3, fork18_outs_2, fork18_outs_1, fork18_outs_0}),
    .outs_valid ({fork18_outs_8_valid, fork18_outs_7_valid, fork18_outs_6_valid, fork18_outs_5_valid, fork18_outs_4_valid, fork18_outs_3_valid, fork18_outs_2_valid, fork18_outs_1_valid, fork18_outs_0_valid}),
    .outs_ready ({fork18_outs_8_ready, fork18_outs_7_ready, fork18_outs_6_ready, fork18_outs_5_ready, fork18_outs_4_ready, fork18_outs_3_ready, fork18_outs_2_ready, fork18_outs_1_ready, fork18_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(36)) cond_br77(
    .condition (fork18_outs_7),
    .condition_valid (fork18_outs_7_valid),
    .condition_ready (fork18_outs_7_ready),
    .data (constant473_outs),
    .data_valid (constant473_outs_valid),
    .data_ready (constant473_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br77_trueOut),
    .trueOut_valid (cond_br77_trueOut_valid),
    .trueOut_ready (cond_br77_trueOut_ready),
    .falseOut (cond_br77_falseOut),
    .falseOut_valid (cond_br77_falseOut_valid),
    .falseOut_ready (cond_br77_falseOut_ready)
  );

  sink #(.DATA_TYPE(36)) sink40(
    .ins (cond_br77_falseOut),
    .ins_valid (cond_br77_falseOut_valid),
    .ins_ready (cond_br77_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(36), .OUTPUT_TYPE(37)) extsi155(
    .ins (cond_br77_trueOut),
    .ins_valid (cond_br77_trueOut_valid),
    .ins_ready (cond_br77_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi155_outs),
    .outs_valid (extsi155_outs_valid),
    .outs_ready (extsi155_outs_ready)
  );

  cond_br #(.DATA_TYPE(33)) cond_br78(
    .condition (fork18_outs_6),
    .condition_valid (fork18_outs_6_valid),
    .condition_ready (fork18_outs_6_ready),
    .data (constant259_outs),
    .data_valid (constant259_outs_valid),
    .data_ready (constant259_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br78_trueOut),
    .trueOut_valid (cond_br78_trueOut_valid),
    .trueOut_ready (cond_br78_trueOut_ready),
    .falseOut (cond_br78_falseOut),
    .falseOut_valid (cond_br78_falseOut_valid),
    .falseOut_ready (cond_br78_falseOut_ready)
  );

  sink #(.DATA_TYPE(33)) sink41(
    .ins (cond_br78_falseOut),
    .ins_valid (cond_br78_falseOut_valid),
    .ins_ready (cond_br78_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br79(
    .condition (fork18_outs_5),
    .condition_valid (fork18_outs_5_valid),
    .condition_ready (fork18_outs_5_ready),
    .data (constant260_outs),
    .data_valid (constant260_outs_valid),
    .data_ready (constant260_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br79_trueOut),
    .trueOut_valid (cond_br79_trueOut_valid),
    .trueOut_ready (cond_br79_trueOut_ready),
    .falseOut (cond_br79_falseOut),
    .falseOut_valid (cond_br79_falseOut_valid),
    .falseOut_ready (cond_br79_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink42(
    .ins (cond_br79_falseOut),
    .ins_valid (cond_br79_falseOut_valid),
    .ins_ready (cond_br79_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(22)) cond_br80(
    .condition (fork18_outs_4),
    .condition_valid (fork18_outs_4_valid),
    .condition_ready (fork18_outs_4_ready),
    .data (constant261_outs),
    .data_valid (constant261_outs_valid),
    .data_ready (constant261_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br80_trueOut),
    .trueOut_valid (cond_br80_trueOut_valid),
    .trueOut_ready (cond_br80_trueOut_ready),
    .falseOut (cond_br80_falseOut),
    .falseOut_valid (cond_br80_falseOut_valid),
    .falseOut_ready (cond_br80_falseOut_ready)
  );

  sink #(.DATA_TYPE(22)) sink43(
    .ins (cond_br80_falseOut),
    .ins_valid (cond_br80_falseOut_valid),
    .ins_ready (cond_br80_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(17)) cond_br81(
    .condition (fork18_outs_3),
    .condition_valid (fork18_outs_3_valid),
    .condition_ready (fork18_outs_3_ready),
    .data (constant262_outs),
    .data_valid (constant262_outs_valid),
    .data_ready (constant262_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br81_trueOut),
    .trueOut_valid (cond_br81_trueOut_valid),
    .trueOut_ready (cond_br81_trueOut_ready),
    .falseOut (cond_br81_falseOut),
    .falseOut_valid (cond_br81_falseOut_valid),
    .falseOut_ready (cond_br81_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink44(
    .ins (cond_br81_falseOut),
    .ins_valid (cond_br81_falseOut_valid),
    .ins_ready (cond_br81_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br82(
    .condition (fork18_outs_2),
    .condition_valid (fork18_outs_2_valid),
    .condition_ready (fork18_outs_2_ready),
    .data (constant263_outs),
    .data_valid (constant263_outs_valid),
    .data_ready (constant263_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br82_trueOut),
    .trueOut_valid (cond_br82_trueOut_valid),
    .trueOut_ready (cond_br82_trueOut_ready),
    .falseOut (cond_br82_falseOut),
    .falseOut_valid (cond_br82_falseOut_valid),
    .falseOut_ready (cond_br82_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink45(
    .ins (cond_br82_falseOut),
    .ins_valid (cond_br82_falseOut_valid),
    .ins_ready (cond_br82_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer24(
    .ins (cond_br74_falseOut),
    .ins_valid (cond_br74_falseOut_valid),
    .ins_ready (cond_br74_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer24_outs),
    .outs_valid (buffer24_outs_valid),
    .outs_ready (buffer24_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer25(
    .ins (buffer24_outs),
    .ins_valid (buffer24_outs_valid),
    .ins_ready (buffer24_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer25_outs),
    .outs_valid (buffer25_outs_valid),
    .outs_ready (buffer25_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br83(
    .condition (fork18_outs_0),
    .condition_valid (fork18_outs_0_valid),
    .condition_ready (fork18_outs_0_ready),
    .data (buffer25_outs),
    .data_valid (buffer25_outs_valid),
    .data_ready (buffer25_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br83_trueOut),
    .trueOut_valid (cond_br83_trueOut_valid),
    .trueOut_ready (cond_br83_trueOut_ready),
    .falseOut (cond_br83_falseOut),
    .falseOut_valid (cond_br83_falseOut_valid),
    .falseOut_ready (cond_br83_falseOut_ready)
  );

  cond_br_dataless cond_br84(
    .condition (fork18_outs_1),
    .condition_valid (fork18_outs_1_valid),
    .condition_ready (fork18_outs_1_ready),
    .data_valid (fork17_outs_6_valid),
    .data_ready (fork17_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br84_trueOut_valid),
    .trueOut_ready (cond_br84_trueOut_ready),
    .falseOut_valid (cond_br84_falseOut_valid),
    .falseOut_ready (cond_br84_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br85(
    .condition (fork18_outs_8),
    .condition_valid (fork18_outs_8_valid),
    .condition_ready (fork18_outs_8_ready),
    .data (fork16_outs_1),
    .data_valid (fork16_outs_1_valid),
    .data_ready (fork16_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br85_trueOut),
    .trueOut_valid (cond_br85_trueOut_valid),
    .trueOut_ready (cond_br85_trueOut_ready),
    .falseOut (cond_br85_falseOut),
    .falseOut_valid (cond_br85_falseOut_valid),
    .falseOut_ready (cond_br85_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink46(
    .ins (cond_br85_trueOut),
    .ins_valid (cond_br85_trueOut_valid),
    .ins_ready (cond_br85_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer32(
    .ins (cond_br85_falseOut),
    .ins_valid (cond_br85_falseOut_valid),
    .ins_ready (cond_br85_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer32_outs),
    .outs_valid (buffer32_outs_valid),
    .outs_ready (buffer32_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer33(
    .ins (buffer32_outs),
    .ins_valid (buffer32_outs_valid),
    .ins_ready (buffer32_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer33_outs),
    .outs_valid (buffer33_outs_valid),
    .outs_ready (buffer33_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork19(
    .ins (buffer33_outs),
    .ins_valid (buffer33_outs_valid),
    .ins_ready (buffer33_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork19_outs_1, fork19_outs_0}),
    .outs_valid ({fork19_outs_1_valid, fork19_outs_0_valid}),
    .outs_ready ({fork19_outs_1_ready, fork19_outs_0_ready})
  );

  oehb_dataless buffer34(
    .ins_valid (cond_br84_falseOut_valid),
    .ins_ready (cond_br84_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer34_outs_valid),
    .outs_ready (buffer34_outs_ready)
  );

  tehb_dataless buffer35(
    .ins_valid (buffer34_outs_valid),
    .ins_ready (buffer34_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer35_outs_valid),
    .outs_ready (buffer35_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork20(
    .ins_valid (buffer35_outs_valid),
    .ins_ready (buffer35_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork20_outs_6_valid, fork20_outs_5_valid, fork20_outs_4_valid, fork20_outs_3_valid, fork20_outs_2_valid, fork20_outs_1_valid, fork20_outs_0_valid}),
    .outs_ready ({fork20_outs_6_ready, fork20_outs_5_ready, fork20_outs_4_ready, fork20_outs_3_ready, fork20_outs_2_ready, fork20_outs_1_ready, fork20_outs_0_ready})
  );

  handshake_constant_43 #(.DATA_WIDTH(36)) constant475(
    .ctrl_valid (fork20_outs_1_valid),
    .ctrl_ready (fork20_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant475_outs),
    .outs_valid (constant475_outs_valid),
    .outs_ready (constant475_outs_ready)
  );

  handshake_constant_44 #(.DATA_WIDTH(32)) constant476(
    .ctrl_valid (fork20_outs_0_valid),
    .ctrl_ready (fork20_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant476_outs),
    .outs_valid (constant476_outs_valid),
    .outs_ready (constant476_outs_ready)
  );

  handshake_constant_45 #(.DATA_WIDTH(27)) constant267(
    .ctrl_valid (fork20_outs_5_valid),
    .ctrl_ready (fork20_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant267_outs),
    .outs_valid (constant267_outs_valid),
    .outs_ready (constant267_outs_ready)
  );

  handshake_constant_46 #(.DATA_WIDTH(22)) constant268(
    .ctrl_valid (fork20_outs_4_valid),
    .ctrl_ready (fork20_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant268_outs),
    .outs_valid (constant268_outs_valid),
    .outs_ready (constant268_outs_ready)
  );

  handshake_constant_47 #(.DATA_WIDTH(17)) constant269(
    .ctrl_valid (fork20_outs_3_valid),
    .ctrl_ready (fork20_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant269_outs),
    .outs_valid (constant269_outs_valid),
    .outs_ready (constant269_outs_ready)
  );

  handshake_constant_48 #(.DATA_WIDTH(12)) constant270(
    .ctrl_valid (fork20_outs_2_valid),
    .ctrl_ready (fork20_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant270_outs),
    .outs_valid (constant270_outs_valid),
    .outs_ready (constant270_outs_ready)
  );

  source source7(
    .clk (clk),
    .rst (rst),
    .outs_valid (source7_outs_valid),
    .outs_ready (source7_outs_ready)
  );

  handshake_constant_49 #(.DATA_WIDTH(4)) constant477(
    .ctrl_valid (source7_outs_valid),
    .ctrl_ready (source7_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant477_outs),
    .outs_valid (constant477_outs_valid),
    .outs_ready (constant477_outs_ready)
  );

  extsi #(.INPUT_TYPE(4), .OUTPUT_TYPE(5)) extsi156(
    .ins (constant477_outs),
    .ins_valid (constant477_outs_valid),
    .ins_ready (constant477_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi156_outs),
    .outs_valid (extsi156_outs_valid),
    .outs_ready (extsi156_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi6(
    .lhs (fork19_outs_0),
    .lhs_valid (fork19_outs_0_valid),
    .lhs_ready (fork19_outs_0_ready),
    .rhs (extsi156_outs),
    .rhs_valid (extsi156_outs_valid),
    .rhs_ready (extsi156_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi6_result),
    .result_valid (cmpi6_result_valid),
    .result_ready (cmpi6_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork21(
    .ins (cmpi6_result),
    .ins_valid (cmpi6_result_valid),
    .ins_ready (cmpi6_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork21_outs_8, fork21_outs_7, fork21_outs_6, fork21_outs_5, fork21_outs_4, fork21_outs_3, fork21_outs_2, fork21_outs_1, fork21_outs_0}),
    .outs_valid ({fork21_outs_8_valid, fork21_outs_7_valid, fork21_outs_6_valid, fork21_outs_5_valid, fork21_outs_4_valid, fork21_outs_3_valid, fork21_outs_2_valid, fork21_outs_1_valid, fork21_outs_0_valid}),
    .outs_ready ({fork21_outs_8_ready, fork21_outs_7_ready, fork21_outs_6_ready, fork21_outs_5_ready, fork21_outs_4_ready, fork21_outs_3_ready, fork21_outs_2_ready, fork21_outs_1_ready, fork21_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(36)) cond_br86(
    .condition (fork21_outs_7),
    .condition_valid (fork21_outs_7_valid),
    .condition_ready (fork21_outs_7_ready),
    .data (constant475_outs),
    .data_valid (constant475_outs_valid),
    .data_ready (constant475_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br86_trueOut),
    .trueOut_valid (cond_br86_trueOut_valid),
    .trueOut_ready (cond_br86_trueOut_ready),
    .falseOut (cond_br86_falseOut),
    .falseOut_valid (cond_br86_falseOut_valid),
    .falseOut_ready (cond_br86_falseOut_ready)
  );

  sink #(.DATA_TYPE(36)) sink48(
    .ins (cond_br86_falseOut),
    .ins_valid (cond_br86_falseOut_valid),
    .ins_ready (cond_br86_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(36), .OUTPUT_TYPE(37)) extsi157(
    .ins (cond_br86_trueOut),
    .ins_valid (cond_br86_trueOut_valid),
    .ins_ready (cond_br86_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi157_outs),
    .outs_valid (extsi157_outs_valid),
    .outs_ready (extsi157_outs_ready)
  );

  cond_br #(.DATA_TYPE(32)) cond_br87(
    .condition (fork21_outs_6),
    .condition_valid (fork21_outs_6_valid),
    .condition_ready (fork21_outs_6_ready),
    .data (constant476_outs),
    .data_valid (constant476_outs_valid),
    .data_ready (constant476_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br87_trueOut),
    .trueOut_valid (cond_br87_trueOut_valid),
    .trueOut_ready (cond_br87_trueOut_ready),
    .falseOut (cond_br87_falseOut),
    .falseOut_valid (cond_br87_falseOut_valid),
    .falseOut_ready (cond_br87_falseOut_ready)
  );

  sink #(.DATA_TYPE(32)) sink49(
    .ins (cond_br87_falseOut),
    .ins_valid (cond_br87_falseOut_valid),
    .ins_ready (cond_br87_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(32), .OUTPUT_TYPE(33)) extsi158(
    .ins (cond_br87_trueOut),
    .ins_valid (cond_br87_trueOut_valid),
    .ins_ready (cond_br87_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi158_outs),
    .outs_valid (extsi158_outs_valid),
    .outs_ready (extsi158_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br88(
    .condition (fork21_outs_5),
    .condition_valid (fork21_outs_5_valid),
    .condition_ready (fork21_outs_5_ready),
    .data (constant267_outs),
    .data_valid (constant267_outs_valid),
    .data_ready (constant267_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br88_trueOut),
    .trueOut_valid (cond_br88_trueOut_valid),
    .trueOut_ready (cond_br88_trueOut_ready),
    .falseOut (cond_br88_falseOut),
    .falseOut_valid (cond_br88_falseOut_valid),
    .falseOut_ready (cond_br88_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink50(
    .ins (cond_br88_falseOut),
    .ins_valid (cond_br88_falseOut_valid),
    .ins_ready (cond_br88_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(22)) cond_br89(
    .condition (fork21_outs_4),
    .condition_valid (fork21_outs_4_valid),
    .condition_ready (fork21_outs_4_ready),
    .data (constant268_outs),
    .data_valid (constant268_outs_valid),
    .data_ready (constant268_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br89_trueOut),
    .trueOut_valid (cond_br89_trueOut_valid),
    .trueOut_ready (cond_br89_trueOut_ready),
    .falseOut (cond_br89_falseOut),
    .falseOut_valid (cond_br89_falseOut_valid),
    .falseOut_ready (cond_br89_falseOut_ready)
  );

  sink #(.DATA_TYPE(22)) sink51(
    .ins (cond_br89_falseOut),
    .ins_valid (cond_br89_falseOut_valid),
    .ins_ready (cond_br89_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(17)) cond_br90(
    .condition (fork21_outs_3),
    .condition_valid (fork21_outs_3_valid),
    .condition_ready (fork21_outs_3_ready),
    .data (constant269_outs),
    .data_valid (constant269_outs_valid),
    .data_ready (constant269_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br90_trueOut),
    .trueOut_valid (cond_br90_trueOut_valid),
    .trueOut_ready (cond_br90_trueOut_ready),
    .falseOut (cond_br90_falseOut),
    .falseOut_valid (cond_br90_falseOut_valid),
    .falseOut_ready (cond_br90_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink52(
    .ins (cond_br90_falseOut),
    .ins_valid (cond_br90_falseOut_valid),
    .ins_ready (cond_br90_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br91(
    .condition (fork21_outs_2),
    .condition_valid (fork21_outs_2_valid),
    .condition_ready (fork21_outs_2_ready),
    .data (constant270_outs),
    .data_valid (constant270_outs_valid),
    .data_ready (constant270_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br91_trueOut),
    .trueOut_valid (cond_br91_trueOut_valid),
    .trueOut_ready (cond_br91_trueOut_ready),
    .falseOut (cond_br91_falseOut),
    .falseOut_valid (cond_br91_falseOut_valid),
    .falseOut_ready (cond_br91_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink53(
    .ins (cond_br91_falseOut),
    .ins_valid (cond_br91_falseOut_valid),
    .ins_ready (cond_br91_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer30(
    .ins (cond_br83_falseOut),
    .ins_valid (cond_br83_falseOut_valid),
    .ins_ready (cond_br83_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer30_outs),
    .outs_valid (buffer30_outs_valid),
    .outs_ready (buffer30_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer31(
    .ins (buffer30_outs),
    .ins_valid (buffer30_outs_valid),
    .ins_ready (buffer30_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer31_outs),
    .outs_valid (buffer31_outs_valid),
    .outs_ready (buffer31_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br92(
    .condition (fork21_outs_0),
    .condition_valid (fork21_outs_0_valid),
    .condition_ready (fork21_outs_0_ready),
    .data (buffer31_outs),
    .data_valid (buffer31_outs_valid),
    .data_ready (buffer31_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br92_trueOut),
    .trueOut_valid (cond_br92_trueOut_valid),
    .trueOut_ready (cond_br92_trueOut_ready),
    .falseOut (cond_br92_falseOut),
    .falseOut_valid (cond_br92_falseOut_valid),
    .falseOut_ready (cond_br92_falseOut_ready)
  );

  cond_br_dataless cond_br93(
    .condition (fork21_outs_1),
    .condition_valid (fork21_outs_1_valid),
    .condition_ready (fork21_outs_1_ready),
    .data_valid (fork20_outs_6_valid),
    .data_ready (fork20_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br93_trueOut_valid),
    .trueOut_ready (cond_br93_trueOut_ready),
    .falseOut_valid (cond_br93_falseOut_valid),
    .falseOut_ready (cond_br93_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br94(
    .condition (fork21_outs_8),
    .condition_valid (fork21_outs_8_valid),
    .condition_ready (fork21_outs_8_ready),
    .data (fork19_outs_1),
    .data_valid (fork19_outs_1_valid),
    .data_ready (fork19_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br94_trueOut),
    .trueOut_valid (cond_br94_trueOut_valid),
    .trueOut_ready (cond_br94_trueOut_ready),
    .falseOut (cond_br94_falseOut),
    .falseOut_valid (cond_br94_falseOut_valid),
    .falseOut_ready (cond_br94_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink54(
    .ins (cond_br94_trueOut),
    .ins_valid (cond_br94_trueOut_valid),
    .ins_ready (cond_br94_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer38(
    .ins (cond_br94_falseOut),
    .ins_valid (cond_br94_falseOut_valid),
    .ins_ready (cond_br94_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer38_outs),
    .outs_valid (buffer38_outs_valid),
    .outs_ready (buffer38_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer39(
    .ins (buffer38_outs),
    .ins_valid (buffer38_outs_valid),
    .ins_ready (buffer38_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer39_outs),
    .outs_valid (buffer39_outs_valid),
    .outs_ready (buffer39_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork22(
    .ins (buffer39_outs),
    .ins_valid (buffer39_outs_valid),
    .ins_ready (buffer39_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork22_outs_1, fork22_outs_0}),
    .outs_valid ({fork22_outs_1_valid, fork22_outs_0_valid}),
    .outs_ready ({fork22_outs_1_ready, fork22_outs_0_ready})
  );

  oehb_dataless buffer40(
    .ins_valid (cond_br93_falseOut_valid),
    .ins_ready (cond_br93_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer40_outs_valid),
    .outs_ready (buffer40_outs_ready)
  );

  tehb_dataless buffer41(
    .ins_valid (buffer40_outs_valid),
    .ins_ready (buffer40_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer41_outs_valid),
    .outs_ready (buffer41_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork23(
    .ins_valid (buffer41_outs_valid),
    .ins_ready (buffer41_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork23_outs_6_valid, fork23_outs_5_valid, fork23_outs_4_valid, fork23_outs_3_valid, fork23_outs_2_valid, fork23_outs_1_valid, fork23_outs_0_valid}),
    .outs_ready ({fork23_outs_6_ready, fork23_outs_5_ready, fork23_outs_4_ready, fork23_outs_3_ready, fork23_outs_2_ready, fork23_outs_1_ready, fork23_outs_0_ready})
  );

  handshake_constant_50 #(.DATA_WIDTH(37)) constant272(
    .ctrl_valid (fork23_outs_5_valid),
    .ctrl_ready (fork23_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant272_outs),
    .outs_valid (constant272_outs_valid),
    .outs_ready (constant272_outs_ready)
  );

  handshake_constant_51 #(.DATA_WIDTH(32)) constant478(
    .ctrl_valid (fork23_outs_1_valid),
    .ctrl_ready (fork23_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant478_outs),
    .outs_valid (constant478_outs_valid),
    .outs_ready (constant478_outs_ready)
  );

  handshake_constant_52 #(.DATA_WIDTH(27)) constant274(
    .ctrl_valid (fork23_outs_4_valid),
    .ctrl_ready (fork23_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant274_outs),
    .outs_valid (constant274_outs_valid),
    .outs_ready (constant274_outs_ready)
  );

  handshake_constant_53 #(.DATA_WIDTH(19)) constant479(
    .ctrl_valid (fork23_outs_0_valid),
    .ctrl_ready (fork23_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant479_outs),
    .outs_valid (constant479_outs_valid),
    .outs_ready (constant479_outs_ready)
  );

  handshake_constant_54 #(.DATA_WIDTH(17)) constant276(
    .ctrl_valid (fork23_outs_3_valid),
    .ctrl_ready (fork23_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant276_outs),
    .outs_valid (constant276_outs_valid),
    .outs_ready (constant276_outs_ready)
  );

  handshake_constant_55 #(.DATA_WIDTH(12)) constant277(
    .ctrl_valid (fork23_outs_2_valid),
    .ctrl_ready (fork23_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant277_outs),
    .outs_valid (constant277_outs_valid),
    .outs_ready (constant277_outs_ready)
  );

  source source8(
    .clk (clk),
    .rst (rst),
    .outs_valid (source8_outs_valid),
    .outs_ready (source8_outs_ready)
  );

  handshake_constant_56 #(.DATA_WIDTH(4)) constant480(
    .ctrl_valid (source8_outs_valid),
    .ctrl_ready (source8_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant480_outs),
    .outs_valid (constant480_outs_valid),
    .outs_ready (constant480_outs_ready)
  );

  extsi #(.INPUT_TYPE(4), .OUTPUT_TYPE(5)) extsi159(
    .ins (constant480_outs),
    .ins_valid (constant480_outs_valid),
    .ins_ready (constant480_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi159_outs),
    .outs_valid (extsi159_outs_valid),
    .outs_ready (extsi159_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi7(
    .lhs (fork22_outs_0),
    .lhs_valid (fork22_outs_0_valid),
    .lhs_ready (fork22_outs_0_ready),
    .rhs (extsi159_outs),
    .rhs_valid (extsi159_outs_valid),
    .rhs_ready (extsi159_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi7_result),
    .result_valid (cmpi7_result_valid),
    .result_ready (cmpi7_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork24(
    .ins (cmpi7_result),
    .ins_valid (cmpi7_result_valid),
    .ins_ready (cmpi7_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork24_outs_8, fork24_outs_7, fork24_outs_6, fork24_outs_5, fork24_outs_4, fork24_outs_3, fork24_outs_2, fork24_outs_1, fork24_outs_0}),
    .outs_valid ({fork24_outs_8_valid, fork24_outs_7_valid, fork24_outs_6_valid, fork24_outs_5_valid, fork24_outs_4_valid, fork24_outs_3_valid, fork24_outs_2_valid, fork24_outs_1_valid, fork24_outs_0_valid}),
    .outs_ready ({fork24_outs_8_ready, fork24_outs_7_ready, fork24_outs_6_ready, fork24_outs_5_ready, fork24_outs_4_ready, fork24_outs_3_ready, fork24_outs_2_ready, fork24_outs_1_ready, fork24_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br95(
    .condition (fork24_outs_5),
    .condition_valid (fork24_outs_5_valid),
    .condition_ready (fork24_outs_5_ready),
    .data (constant272_outs),
    .data_valid (constant272_outs_valid),
    .data_ready (constant272_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br95_trueOut),
    .trueOut_valid (cond_br95_trueOut_valid),
    .trueOut_ready (cond_br95_trueOut_ready),
    .falseOut (cond_br95_falseOut),
    .falseOut_valid (cond_br95_falseOut_valid),
    .falseOut_ready (cond_br95_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink56(
    .ins (cond_br95_falseOut),
    .ins_valid (cond_br95_falseOut_valid),
    .ins_ready (cond_br95_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(32)) cond_br96(
    .condition (fork24_outs_7),
    .condition_valid (fork24_outs_7_valid),
    .condition_ready (fork24_outs_7_ready),
    .data (constant478_outs),
    .data_valid (constant478_outs_valid),
    .data_ready (constant478_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br96_trueOut),
    .trueOut_valid (cond_br96_trueOut_valid),
    .trueOut_ready (cond_br96_trueOut_ready),
    .falseOut (cond_br96_falseOut),
    .falseOut_valid (cond_br96_falseOut_valid),
    .falseOut_ready (cond_br96_falseOut_ready)
  );

  sink #(.DATA_TYPE(32)) sink57(
    .ins (cond_br96_falseOut),
    .ins_valid (cond_br96_falseOut_valid),
    .ins_ready (cond_br96_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(32), .OUTPUT_TYPE(33)) extsi160(
    .ins (cond_br96_trueOut),
    .ins_valid (cond_br96_trueOut_valid),
    .ins_ready (cond_br96_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi160_outs),
    .outs_valid (extsi160_outs_valid),
    .outs_ready (extsi160_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br97(
    .condition (fork24_outs_4),
    .condition_valid (fork24_outs_4_valid),
    .condition_ready (fork24_outs_4_ready),
    .data (constant274_outs),
    .data_valid (constant274_outs_valid),
    .data_ready (constant274_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br97_trueOut),
    .trueOut_valid (cond_br97_trueOut_valid),
    .trueOut_ready (cond_br97_trueOut_ready),
    .falseOut (cond_br97_falseOut),
    .falseOut_valid (cond_br97_falseOut_valid),
    .falseOut_ready (cond_br97_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink58(
    .ins (cond_br97_falseOut),
    .ins_valid (cond_br97_falseOut_valid),
    .ins_ready (cond_br97_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(19)) cond_br98(
    .condition (fork24_outs_6),
    .condition_valid (fork24_outs_6_valid),
    .condition_ready (fork24_outs_6_ready),
    .data (constant479_outs),
    .data_valid (constant479_outs_valid),
    .data_ready (constant479_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br98_trueOut),
    .trueOut_valid (cond_br98_trueOut_valid),
    .trueOut_ready (cond_br98_trueOut_ready),
    .falseOut (cond_br98_falseOut),
    .falseOut_valid (cond_br98_falseOut_valid),
    .falseOut_ready (cond_br98_falseOut_ready)
  );

  sink #(.DATA_TYPE(19)) sink59(
    .ins (cond_br98_falseOut),
    .ins_valid (cond_br98_falseOut_valid),
    .ins_ready (cond_br98_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(19), .OUTPUT_TYPE(22)) extsi161(
    .ins (cond_br98_trueOut),
    .ins_valid (cond_br98_trueOut_valid),
    .ins_ready (cond_br98_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi161_outs),
    .outs_valid (extsi161_outs_valid),
    .outs_ready (extsi161_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br99(
    .condition (fork24_outs_3),
    .condition_valid (fork24_outs_3_valid),
    .condition_ready (fork24_outs_3_ready),
    .data (constant276_outs),
    .data_valid (constant276_outs_valid),
    .data_ready (constant276_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br99_trueOut),
    .trueOut_valid (cond_br99_trueOut_valid),
    .trueOut_ready (cond_br99_trueOut_ready),
    .falseOut (cond_br99_falseOut),
    .falseOut_valid (cond_br99_falseOut_valid),
    .falseOut_ready (cond_br99_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink60(
    .ins (cond_br99_falseOut),
    .ins_valid (cond_br99_falseOut_valid),
    .ins_ready (cond_br99_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br100(
    .condition (fork24_outs_2),
    .condition_valid (fork24_outs_2_valid),
    .condition_ready (fork24_outs_2_ready),
    .data (constant277_outs),
    .data_valid (constant277_outs_valid),
    .data_ready (constant277_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br100_trueOut),
    .trueOut_valid (cond_br100_trueOut_valid),
    .trueOut_ready (cond_br100_trueOut_ready),
    .falseOut (cond_br100_falseOut),
    .falseOut_valid (cond_br100_falseOut_valid),
    .falseOut_ready (cond_br100_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink61(
    .ins (cond_br100_falseOut),
    .ins_valid (cond_br100_falseOut_valid),
    .ins_ready (cond_br100_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer36(
    .ins (cond_br92_falseOut),
    .ins_valid (cond_br92_falseOut_valid),
    .ins_ready (cond_br92_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer36_outs),
    .outs_valid (buffer36_outs_valid),
    .outs_ready (buffer36_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer37(
    .ins (buffer36_outs),
    .ins_valid (buffer36_outs_valid),
    .ins_ready (buffer36_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer37_outs),
    .outs_valid (buffer37_outs_valid),
    .outs_ready (buffer37_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br101(
    .condition (fork24_outs_0),
    .condition_valid (fork24_outs_0_valid),
    .condition_ready (fork24_outs_0_ready),
    .data (buffer37_outs),
    .data_valid (buffer37_outs_valid),
    .data_ready (buffer37_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br101_trueOut),
    .trueOut_valid (cond_br101_trueOut_valid),
    .trueOut_ready (cond_br101_trueOut_ready),
    .falseOut (cond_br101_falseOut),
    .falseOut_valid (cond_br101_falseOut_valid),
    .falseOut_ready (cond_br101_falseOut_ready)
  );

  cond_br_dataless cond_br102(
    .condition (fork24_outs_1),
    .condition_valid (fork24_outs_1_valid),
    .condition_ready (fork24_outs_1_ready),
    .data_valid (fork23_outs_6_valid),
    .data_ready (fork23_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br102_trueOut_valid),
    .trueOut_ready (cond_br102_trueOut_ready),
    .falseOut_valid (cond_br102_falseOut_valid),
    .falseOut_ready (cond_br102_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br103(
    .condition (fork24_outs_8),
    .condition_valid (fork24_outs_8_valid),
    .condition_ready (fork24_outs_8_ready),
    .data (fork22_outs_1),
    .data_valid (fork22_outs_1_valid),
    .data_ready (fork22_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br103_trueOut),
    .trueOut_valid (cond_br103_trueOut_valid),
    .trueOut_ready (cond_br103_trueOut_ready),
    .falseOut (cond_br103_falseOut),
    .falseOut_valid (cond_br103_falseOut_valid),
    .falseOut_ready (cond_br103_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink62(
    .ins (cond_br103_trueOut),
    .ins_valid (cond_br103_trueOut_valid),
    .ins_ready (cond_br103_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer44(
    .ins (cond_br103_falseOut),
    .ins_valid (cond_br103_falseOut_valid),
    .ins_ready (cond_br103_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer44_outs),
    .outs_valid (buffer44_outs_valid),
    .outs_ready (buffer44_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer45(
    .ins (buffer44_outs),
    .ins_valid (buffer44_outs_valid),
    .ins_ready (buffer44_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer45_outs),
    .outs_valid (buffer45_outs_valid),
    .outs_ready (buffer45_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork25(
    .ins (buffer45_outs),
    .ins_valid (buffer45_outs_valid),
    .ins_ready (buffer45_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork25_outs_1, fork25_outs_0}),
    .outs_valid ({fork25_outs_1_valid, fork25_outs_0_valid}),
    .outs_ready ({fork25_outs_1_ready, fork25_outs_0_ready})
  );

  oehb_dataless buffer46(
    .ins_valid (cond_br102_falseOut_valid),
    .ins_ready (cond_br102_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer46_outs_valid),
    .outs_ready (buffer46_outs_ready)
  );

  tehb_dataless buffer47(
    .ins_valid (buffer46_outs_valid),
    .ins_ready (buffer46_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer47_outs_valid),
    .outs_ready (buffer47_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork26(
    .ins_valid (buffer47_outs_valid),
    .ins_ready (buffer47_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork26_outs_6_valid, fork26_outs_5_valid, fork26_outs_4_valid, fork26_outs_3_valid, fork26_outs_2_valid, fork26_outs_1_valid, fork26_outs_0_valid}),
    .outs_ready ({fork26_outs_6_ready, fork26_outs_5_ready, fork26_outs_4_ready, fork26_outs_3_ready, fork26_outs_2_ready, fork26_outs_1_ready, fork26_outs_0_ready})
  );

  handshake_constant_57 #(.DATA_WIDTH(37)) constant279(
    .ctrl_valid (fork26_outs_5_valid),
    .ctrl_ready (fork26_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant279_outs),
    .outs_valid (constant279_outs_valid),
    .outs_ready (constant279_outs_ready)
  );

  handshake_constant_58 #(.DATA_WIDTH(32)) constant481(
    .ctrl_valid (fork26_outs_2_valid),
    .ctrl_ready (fork26_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant481_outs),
    .outs_valid (constant481_outs_valid),
    .outs_ready (constant481_outs_ready)
  );

  handshake_constant_59 #(.DATA_WIDTH(27)) constant281(
    .ctrl_valid (fork26_outs_4_valid),
    .ctrl_ready (fork26_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant281_outs),
    .outs_valid (constant281_outs_valid),
    .outs_ready (constant281_outs_ready)
  );

  handshake_constant_60 #(.DATA_WIDTH(20)) constant482(
    .ctrl_valid (fork26_outs_1_valid),
    .ctrl_ready (fork26_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant482_outs),
    .outs_valid (constant482_outs_valid),
    .outs_ready (constant482_outs_ready)
  );

  handshake_constant_61 #(.DATA_WIDTH(16)) constant483(
    .ctrl_valid (fork26_outs_0_valid),
    .ctrl_ready (fork26_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant483_outs),
    .outs_valid (constant483_outs_valid),
    .outs_ready (constant483_outs_ready)
  );

  handshake_constant_62 #(.DATA_WIDTH(12)) constant284(
    .ctrl_valid (fork26_outs_3_valid),
    .ctrl_ready (fork26_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant284_outs),
    .outs_valid (constant284_outs_valid),
    .outs_ready (constant284_outs_ready)
  );

  source source9(
    .clk (clk),
    .rst (rst),
    .outs_valid (source9_outs_valid),
    .outs_ready (source9_outs_ready)
  );

  handshake_constant_63 #(.DATA_WIDTH(5)) constant484(
    .ctrl_valid (source9_outs_valid),
    .ctrl_ready (source9_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant484_outs),
    .outs_valid (constant484_outs_valid),
    .outs_ready (constant484_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi8(
    .lhs (fork25_outs_0),
    .lhs_valid (fork25_outs_0_valid),
    .lhs_ready (fork25_outs_0_ready),
    .rhs (constant484_outs),
    .rhs_valid (constant484_outs_valid),
    .rhs_ready (constant484_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi8_result),
    .result_valid (cmpi8_result_valid),
    .result_ready (cmpi8_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork27(
    .ins (cmpi8_result),
    .ins_valid (cmpi8_result_valid),
    .ins_ready (cmpi8_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork27_outs_8, fork27_outs_7, fork27_outs_6, fork27_outs_5, fork27_outs_4, fork27_outs_3, fork27_outs_2, fork27_outs_1, fork27_outs_0}),
    .outs_valid ({fork27_outs_8_valid, fork27_outs_7_valid, fork27_outs_6_valid, fork27_outs_5_valid, fork27_outs_4_valid, fork27_outs_3_valid, fork27_outs_2_valid, fork27_outs_1_valid, fork27_outs_0_valid}),
    .outs_ready ({fork27_outs_8_ready, fork27_outs_7_ready, fork27_outs_6_ready, fork27_outs_5_ready, fork27_outs_4_ready, fork27_outs_3_ready, fork27_outs_2_ready, fork27_outs_1_ready, fork27_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br104(
    .condition (fork27_outs_4),
    .condition_valid (fork27_outs_4_valid),
    .condition_ready (fork27_outs_4_ready),
    .data (constant279_outs),
    .data_valid (constant279_outs_valid),
    .data_ready (constant279_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br104_trueOut),
    .trueOut_valid (cond_br104_trueOut_valid),
    .trueOut_ready (cond_br104_trueOut_ready),
    .falseOut (cond_br104_falseOut),
    .falseOut_valid (cond_br104_falseOut_valid),
    .falseOut_ready (cond_br104_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink64(
    .ins (cond_br104_falseOut),
    .ins_valid (cond_br104_falseOut_valid),
    .ins_ready (cond_br104_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(32)) cond_br105(
    .condition (fork27_outs_7),
    .condition_valid (fork27_outs_7_valid),
    .condition_ready (fork27_outs_7_ready),
    .data (constant481_outs),
    .data_valid (constant481_outs_valid),
    .data_ready (constant481_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br105_trueOut),
    .trueOut_valid (cond_br105_trueOut_valid),
    .trueOut_ready (cond_br105_trueOut_ready),
    .falseOut (cond_br105_falseOut),
    .falseOut_valid (cond_br105_falseOut_valid),
    .falseOut_ready (cond_br105_falseOut_ready)
  );

  sink #(.DATA_TYPE(32)) sink65(
    .ins (cond_br105_falseOut),
    .ins_valid (cond_br105_falseOut_valid),
    .ins_ready (cond_br105_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(32), .OUTPUT_TYPE(33)) extsi162(
    .ins (cond_br105_trueOut),
    .ins_valid (cond_br105_trueOut_valid),
    .ins_ready (cond_br105_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi162_outs),
    .outs_valid (extsi162_outs_valid),
    .outs_ready (extsi162_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br106(
    .condition (fork27_outs_3),
    .condition_valid (fork27_outs_3_valid),
    .condition_ready (fork27_outs_3_ready),
    .data (constant281_outs),
    .data_valid (constant281_outs_valid),
    .data_ready (constant281_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br106_trueOut),
    .trueOut_valid (cond_br106_trueOut_valid),
    .trueOut_ready (cond_br106_trueOut_ready),
    .falseOut (cond_br106_falseOut),
    .falseOut_valid (cond_br106_falseOut_valid),
    .falseOut_ready (cond_br106_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink66(
    .ins (cond_br106_falseOut),
    .ins_valid (cond_br106_falseOut_valid),
    .ins_ready (cond_br106_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(20)) cond_br107(
    .condition (fork27_outs_6),
    .condition_valid (fork27_outs_6_valid),
    .condition_ready (fork27_outs_6_ready),
    .data (constant482_outs),
    .data_valid (constant482_outs_valid),
    .data_ready (constant482_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br107_trueOut),
    .trueOut_valid (cond_br107_trueOut_valid),
    .trueOut_ready (cond_br107_trueOut_ready),
    .falseOut (cond_br107_falseOut),
    .falseOut_valid (cond_br107_falseOut_valid),
    .falseOut_ready (cond_br107_falseOut_ready)
  );

  sink #(.DATA_TYPE(20)) sink67(
    .ins (cond_br107_falseOut),
    .ins_valid (cond_br107_falseOut_valid),
    .ins_ready (cond_br107_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(20), .OUTPUT_TYPE(22)) extsi163(
    .ins (cond_br107_trueOut),
    .ins_valid (cond_br107_trueOut_valid),
    .ins_ready (cond_br107_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi163_outs),
    .outs_valid (extsi163_outs_valid),
    .outs_ready (extsi163_outs_ready)
  );

  cond_br #(.DATA_TYPE(16)) cond_br108(
    .condition (fork27_outs_5),
    .condition_valid (fork27_outs_5_valid),
    .condition_ready (fork27_outs_5_ready),
    .data (constant483_outs),
    .data_valid (constant483_outs_valid),
    .data_ready (constant483_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br108_trueOut),
    .trueOut_valid (cond_br108_trueOut_valid),
    .trueOut_ready (cond_br108_trueOut_ready),
    .falseOut (cond_br108_falseOut),
    .falseOut_valid (cond_br108_falseOut_valid),
    .falseOut_ready (cond_br108_falseOut_ready)
  );

  sink #(.DATA_TYPE(16)) sink68(
    .ins (cond_br108_falseOut),
    .ins_valid (cond_br108_falseOut_valid),
    .ins_ready (cond_br108_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(16), .OUTPUT_TYPE(17)) extsi164(
    .ins (cond_br108_trueOut),
    .ins_valid (cond_br108_trueOut_valid),
    .ins_ready (cond_br108_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi164_outs),
    .outs_valid (extsi164_outs_valid),
    .outs_ready (extsi164_outs_ready)
  );

  cond_br #(.DATA_TYPE(12)) cond_br109(
    .condition (fork27_outs_2),
    .condition_valid (fork27_outs_2_valid),
    .condition_ready (fork27_outs_2_ready),
    .data (constant284_outs),
    .data_valid (constant284_outs_valid),
    .data_ready (constant284_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br109_trueOut),
    .trueOut_valid (cond_br109_trueOut_valid),
    .trueOut_ready (cond_br109_trueOut_ready),
    .falseOut (cond_br109_falseOut),
    .falseOut_valid (cond_br109_falseOut_valid),
    .falseOut_ready (cond_br109_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink69(
    .ins (cond_br109_falseOut),
    .ins_valid (cond_br109_falseOut_valid),
    .ins_ready (cond_br109_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer42(
    .ins (cond_br101_falseOut),
    .ins_valid (cond_br101_falseOut_valid),
    .ins_ready (cond_br101_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer42_outs),
    .outs_valid (buffer42_outs_valid),
    .outs_ready (buffer42_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer43(
    .ins (buffer42_outs),
    .ins_valid (buffer42_outs_valid),
    .ins_ready (buffer42_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer43_outs),
    .outs_valid (buffer43_outs_valid),
    .outs_ready (buffer43_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br110(
    .condition (fork27_outs_0),
    .condition_valid (fork27_outs_0_valid),
    .condition_ready (fork27_outs_0_ready),
    .data (buffer43_outs),
    .data_valid (buffer43_outs_valid),
    .data_ready (buffer43_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br110_trueOut),
    .trueOut_valid (cond_br110_trueOut_valid),
    .trueOut_ready (cond_br110_trueOut_ready),
    .falseOut (cond_br110_falseOut),
    .falseOut_valid (cond_br110_falseOut_valid),
    .falseOut_ready (cond_br110_falseOut_ready)
  );

  cond_br_dataless cond_br111(
    .condition (fork27_outs_1),
    .condition_valid (fork27_outs_1_valid),
    .condition_ready (fork27_outs_1_ready),
    .data_valid (fork26_outs_6_valid),
    .data_ready (fork26_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br111_trueOut_valid),
    .trueOut_ready (cond_br111_trueOut_ready),
    .falseOut_valid (cond_br111_falseOut_valid),
    .falseOut_ready (cond_br111_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br112(
    .condition (fork27_outs_8),
    .condition_valid (fork27_outs_8_valid),
    .condition_ready (fork27_outs_8_ready),
    .data (fork25_outs_1),
    .data_valid (fork25_outs_1_valid),
    .data_ready (fork25_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br112_trueOut),
    .trueOut_valid (cond_br112_trueOut_valid),
    .trueOut_ready (cond_br112_trueOut_ready),
    .falseOut (cond_br112_falseOut),
    .falseOut_valid (cond_br112_falseOut_valid),
    .falseOut_ready (cond_br112_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink70(
    .ins (cond_br112_trueOut),
    .ins_valid (cond_br112_trueOut_valid),
    .ins_ready (cond_br112_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer50(
    .ins (cond_br112_falseOut),
    .ins_valid (cond_br112_falseOut_valid),
    .ins_ready (cond_br112_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer50_outs),
    .outs_valid (buffer50_outs_valid),
    .outs_ready (buffer50_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer51(
    .ins (buffer50_outs),
    .ins_valid (buffer50_outs_valid),
    .ins_ready (buffer50_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer51_outs),
    .outs_valid (buffer51_outs_valid),
    .outs_ready (buffer51_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork28(
    .ins (buffer51_outs),
    .ins_valid (buffer51_outs_valid),
    .ins_ready (buffer51_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork28_outs_1, fork28_outs_0}),
    .outs_valid ({fork28_outs_1_valid, fork28_outs_0_valid}),
    .outs_ready ({fork28_outs_1_ready, fork28_outs_0_ready})
  );

  oehb_dataless buffer52(
    .ins_valid (cond_br111_falseOut_valid),
    .ins_ready (cond_br111_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer52_outs_valid),
    .outs_ready (buffer52_outs_ready)
  );

  tehb_dataless buffer53(
    .ins_valid (buffer52_outs_valid),
    .ins_ready (buffer52_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer53_outs_valid),
    .outs_ready (buffer53_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork29(
    .ins_valid (buffer53_outs_valid),
    .ins_ready (buffer53_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork29_outs_6_valid, fork29_outs_5_valid, fork29_outs_4_valid, fork29_outs_3_valid, fork29_outs_2_valid, fork29_outs_1_valid, fork29_outs_0_valid}),
    .outs_ready ({fork29_outs_6_ready, fork29_outs_5_ready, fork29_outs_4_ready, fork29_outs_3_ready, fork29_outs_2_ready, fork29_outs_1_ready, fork29_outs_0_ready})
  );

  handshake_constant_64 #(.DATA_WIDTH(37)) constant286(
    .ctrl_valid (fork29_outs_5_valid),
    .ctrl_ready (fork29_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant286_outs),
    .outs_valid (constant286_outs_valid),
    .outs_ready (constant286_outs_ready)
  );

  handshake_constant_65 #(.DATA_WIDTH(32)) constant485(
    .ctrl_valid (fork29_outs_2_valid),
    .ctrl_ready (fork29_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant485_outs),
    .outs_valid (constant485_outs_valid),
    .outs_ready (constant485_outs_ready)
  );

  handshake_constant_66 #(.DATA_WIDTH(27)) constant288(
    .ctrl_valid (fork29_outs_4_valid),
    .ctrl_ready (fork29_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant288_outs),
    .outs_valid (constant288_outs_valid),
    .outs_ready (constant288_outs_ready)
  );

  handshake_constant_67 #(.DATA_WIDTH(21)) constant486(
    .ctrl_valid (fork29_outs_1_valid),
    .ctrl_ready (fork29_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant486_outs),
    .outs_valid (constant486_outs_valid),
    .outs_ready (constant486_outs_ready)
  );

  handshake_constant_68 #(.DATA_WIDTH(16)) constant487(
    .ctrl_valid (fork29_outs_0_valid),
    .ctrl_ready (fork29_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant487_outs),
    .outs_valid (constant487_outs_valid),
    .outs_ready (constant487_outs_ready)
  );

  handshake_constant_69 #(.DATA_WIDTH(12)) constant291(
    .ctrl_valid (fork29_outs_3_valid),
    .ctrl_ready (fork29_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant291_outs),
    .outs_valid (constant291_outs_valid),
    .outs_ready (constant291_outs_ready)
  );

  source source10(
    .clk (clk),
    .rst (rst),
    .outs_valid (source10_outs_valid),
    .outs_ready (source10_outs_ready)
  );

  handshake_constant_70 #(.DATA_WIDTH(5)) constant488(
    .ctrl_valid (source10_outs_valid),
    .ctrl_ready (source10_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant488_outs),
    .outs_valid (constant488_outs_valid),
    .outs_ready (constant488_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi9(
    .lhs (fork28_outs_0),
    .lhs_valid (fork28_outs_0_valid),
    .lhs_ready (fork28_outs_0_ready),
    .rhs (constant488_outs),
    .rhs_valid (constant488_outs_valid),
    .rhs_ready (constant488_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi9_result),
    .result_valid (cmpi9_result_valid),
    .result_ready (cmpi9_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork30(
    .ins (cmpi9_result),
    .ins_valid (cmpi9_result_valid),
    .ins_ready (cmpi9_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork30_outs_8, fork30_outs_7, fork30_outs_6, fork30_outs_5, fork30_outs_4, fork30_outs_3, fork30_outs_2, fork30_outs_1, fork30_outs_0}),
    .outs_valid ({fork30_outs_8_valid, fork30_outs_7_valid, fork30_outs_6_valid, fork30_outs_5_valid, fork30_outs_4_valid, fork30_outs_3_valid, fork30_outs_2_valid, fork30_outs_1_valid, fork30_outs_0_valid}),
    .outs_ready ({fork30_outs_8_ready, fork30_outs_7_ready, fork30_outs_6_ready, fork30_outs_5_ready, fork30_outs_4_ready, fork30_outs_3_ready, fork30_outs_2_ready, fork30_outs_1_ready, fork30_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br113(
    .condition (fork30_outs_4),
    .condition_valid (fork30_outs_4_valid),
    .condition_ready (fork30_outs_4_ready),
    .data (constant286_outs),
    .data_valid (constant286_outs_valid),
    .data_ready (constant286_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br113_trueOut),
    .trueOut_valid (cond_br113_trueOut_valid),
    .trueOut_ready (cond_br113_trueOut_ready),
    .falseOut (cond_br113_falseOut),
    .falseOut_valid (cond_br113_falseOut_valid),
    .falseOut_ready (cond_br113_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink72(
    .ins (cond_br113_falseOut),
    .ins_valid (cond_br113_falseOut_valid),
    .ins_ready (cond_br113_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(32)) cond_br114(
    .condition (fork30_outs_7),
    .condition_valid (fork30_outs_7_valid),
    .condition_ready (fork30_outs_7_ready),
    .data (constant485_outs),
    .data_valid (constant485_outs_valid),
    .data_ready (constant485_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br114_trueOut),
    .trueOut_valid (cond_br114_trueOut_valid),
    .trueOut_ready (cond_br114_trueOut_ready),
    .falseOut (cond_br114_falseOut),
    .falseOut_valid (cond_br114_falseOut_valid),
    .falseOut_ready (cond_br114_falseOut_ready)
  );

  sink #(.DATA_TYPE(32)) sink73(
    .ins (cond_br114_falseOut),
    .ins_valid (cond_br114_falseOut_valid),
    .ins_ready (cond_br114_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(32), .OUTPUT_TYPE(33)) extsi165(
    .ins (cond_br114_trueOut),
    .ins_valid (cond_br114_trueOut_valid),
    .ins_ready (cond_br114_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi165_outs),
    .outs_valid (extsi165_outs_valid),
    .outs_ready (extsi165_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br115(
    .condition (fork30_outs_3),
    .condition_valid (fork30_outs_3_valid),
    .condition_ready (fork30_outs_3_ready),
    .data (constant288_outs),
    .data_valid (constant288_outs_valid),
    .data_ready (constant288_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br115_trueOut),
    .trueOut_valid (cond_br115_trueOut_valid),
    .trueOut_ready (cond_br115_trueOut_ready),
    .falseOut (cond_br115_falseOut),
    .falseOut_valid (cond_br115_falseOut_valid),
    .falseOut_ready (cond_br115_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink74(
    .ins (cond_br115_falseOut),
    .ins_valid (cond_br115_falseOut_valid),
    .ins_ready (cond_br115_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(21)) cond_br116(
    .condition (fork30_outs_6),
    .condition_valid (fork30_outs_6_valid),
    .condition_ready (fork30_outs_6_ready),
    .data (constant486_outs),
    .data_valid (constant486_outs_valid),
    .data_ready (constant486_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br116_trueOut),
    .trueOut_valid (cond_br116_trueOut_valid),
    .trueOut_ready (cond_br116_trueOut_ready),
    .falseOut (cond_br116_falseOut),
    .falseOut_valid (cond_br116_falseOut_valid),
    .falseOut_ready (cond_br116_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink75(
    .ins (cond_br116_falseOut),
    .ins_valid (cond_br116_falseOut_valid),
    .ins_ready (cond_br116_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(21), .OUTPUT_TYPE(22)) extsi166(
    .ins (cond_br116_trueOut),
    .ins_valid (cond_br116_trueOut_valid),
    .ins_ready (cond_br116_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi166_outs),
    .outs_valid (extsi166_outs_valid),
    .outs_ready (extsi166_outs_ready)
  );

  cond_br #(.DATA_TYPE(16)) cond_br117(
    .condition (fork30_outs_5),
    .condition_valid (fork30_outs_5_valid),
    .condition_ready (fork30_outs_5_ready),
    .data (constant487_outs),
    .data_valid (constant487_outs_valid),
    .data_ready (constant487_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br117_trueOut),
    .trueOut_valid (cond_br117_trueOut_valid),
    .trueOut_ready (cond_br117_trueOut_ready),
    .falseOut (cond_br117_falseOut),
    .falseOut_valid (cond_br117_falseOut_valid),
    .falseOut_ready (cond_br117_falseOut_ready)
  );

  sink #(.DATA_TYPE(16)) sink76(
    .ins (cond_br117_falseOut),
    .ins_valid (cond_br117_falseOut_valid),
    .ins_ready (cond_br117_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(16), .OUTPUT_TYPE(17)) extsi167(
    .ins (cond_br117_trueOut),
    .ins_valid (cond_br117_trueOut_valid),
    .ins_ready (cond_br117_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi167_outs),
    .outs_valid (extsi167_outs_valid),
    .outs_ready (extsi167_outs_ready)
  );

  cond_br #(.DATA_TYPE(12)) cond_br118(
    .condition (fork30_outs_2),
    .condition_valid (fork30_outs_2_valid),
    .condition_ready (fork30_outs_2_ready),
    .data (constant291_outs),
    .data_valid (constant291_outs_valid),
    .data_ready (constant291_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br118_trueOut),
    .trueOut_valid (cond_br118_trueOut_valid),
    .trueOut_ready (cond_br118_trueOut_ready),
    .falseOut (cond_br118_falseOut),
    .falseOut_valid (cond_br118_falseOut_valid),
    .falseOut_ready (cond_br118_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink77(
    .ins (cond_br118_falseOut),
    .ins_valid (cond_br118_falseOut_valid),
    .ins_ready (cond_br118_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer48(
    .ins (cond_br110_falseOut),
    .ins_valid (cond_br110_falseOut_valid),
    .ins_ready (cond_br110_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer48_outs),
    .outs_valid (buffer48_outs_valid),
    .outs_ready (buffer48_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer49(
    .ins (buffer48_outs),
    .ins_valid (buffer48_outs_valid),
    .ins_ready (buffer48_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer49_outs),
    .outs_valid (buffer49_outs_valid),
    .outs_ready (buffer49_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br119(
    .condition (fork30_outs_0),
    .condition_valid (fork30_outs_0_valid),
    .condition_ready (fork30_outs_0_ready),
    .data (buffer49_outs),
    .data_valid (buffer49_outs_valid),
    .data_ready (buffer49_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br119_trueOut),
    .trueOut_valid (cond_br119_trueOut_valid),
    .trueOut_ready (cond_br119_trueOut_ready),
    .falseOut (cond_br119_falseOut),
    .falseOut_valid (cond_br119_falseOut_valid),
    .falseOut_ready (cond_br119_falseOut_ready)
  );

  cond_br_dataless cond_br120(
    .condition (fork30_outs_1),
    .condition_valid (fork30_outs_1_valid),
    .condition_ready (fork30_outs_1_ready),
    .data_valid (fork29_outs_6_valid),
    .data_ready (fork29_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br120_trueOut_valid),
    .trueOut_ready (cond_br120_trueOut_ready),
    .falseOut_valid (cond_br120_falseOut_valid),
    .falseOut_ready (cond_br120_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br121(
    .condition (fork30_outs_8),
    .condition_valid (fork30_outs_8_valid),
    .condition_ready (fork30_outs_8_ready),
    .data (fork28_outs_1),
    .data_valid (fork28_outs_1_valid),
    .data_ready (fork28_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br121_trueOut),
    .trueOut_valid (cond_br121_trueOut_valid),
    .trueOut_ready (cond_br121_trueOut_ready),
    .falseOut (cond_br121_falseOut),
    .falseOut_valid (cond_br121_falseOut_valid),
    .falseOut_ready (cond_br121_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink78(
    .ins (cond_br121_trueOut),
    .ins_valid (cond_br121_trueOut_valid),
    .ins_ready (cond_br121_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer56(
    .ins (cond_br121_falseOut),
    .ins_valid (cond_br121_falseOut_valid),
    .ins_ready (cond_br121_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer56_outs),
    .outs_valid (buffer56_outs_valid),
    .outs_ready (buffer56_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer57(
    .ins (buffer56_outs),
    .ins_valid (buffer56_outs_valid),
    .ins_ready (buffer56_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer57_outs),
    .outs_valid (buffer57_outs_valid),
    .outs_ready (buffer57_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork31(
    .ins (buffer57_outs),
    .ins_valid (buffer57_outs_valid),
    .ins_ready (buffer57_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork31_outs_1, fork31_outs_0}),
    .outs_valid ({fork31_outs_1_valid, fork31_outs_0_valid}),
    .outs_ready ({fork31_outs_1_ready, fork31_outs_0_ready})
  );

  oehb_dataless buffer58(
    .ins_valid (cond_br120_falseOut_valid),
    .ins_ready (cond_br120_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer58_outs_valid),
    .outs_ready (buffer58_outs_ready)
  );

  tehb_dataless buffer59(
    .ins_valid (buffer58_outs_valid),
    .ins_ready (buffer58_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer59_outs_valid),
    .outs_ready (buffer59_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork32(
    .ins_valid (buffer59_outs_valid),
    .ins_ready (buffer59_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork32_outs_6_valid, fork32_outs_5_valid, fork32_outs_4_valid, fork32_outs_3_valid, fork32_outs_2_valid, fork32_outs_1_valid, fork32_outs_0_valid}),
    .outs_ready ({fork32_outs_6_ready, fork32_outs_5_ready, fork32_outs_4_ready, fork32_outs_3_ready, fork32_outs_2_ready, fork32_outs_1_ready, fork32_outs_0_ready})
  );

  handshake_constant_71 #(.DATA_WIDTH(37)) constant293(
    .ctrl_valid (fork32_outs_5_valid),
    .ctrl_ready (fork32_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant293_outs),
    .outs_valid (constant293_outs_valid),
    .outs_ready (constant293_outs_ready)
  );

  handshake_constant_72 #(.DATA_WIDTH(32)) constant489(
    .ctrl_valid (fork32_outs_2_valid),
    .ctrl_ready (fork32_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant489_outs),
    .outs_valid (constant489_outs_valid),
    .outs_ready (constant489_outs_ready)
  );

  handshake_constant_73 #(.DATA_WIDTH(27)) constant295(
    .ctrl_valid (fork32_outs_4_valid),
    .ctrl_ready (fork32_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant295_outs),
    .outs_valid (constant295_outs_valid),
    .outs_ready (constant295_outs_ready)
  );

  handshake_constant_74 #(.DATA_WIDTH(21)) constant490(
    .ctrl_valid (fork32_outs_1_valid),
    .ctrl_ready (fork32_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant490_outs),
    .outs_valid (constant490_outs_valid),
    .outs_ready (constant490_outs_ready)
  );

  handshake_constant_75 #(.DATA_WIDTH(15)) constant491(
    .ctrl_valid (fork32_outs_0_valid),
    .ctrl_ready (fork32_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant491_outs),
    .outs_valid (constant491_outs_valid),
    .outs_ready (constant491_outs_ready)
  );

  handshake_constant_76 #(.DATA_WIDTH(12)) constant298(
    .ctrl_valid (fork32_outs_3_valid),
    .ctrl_ready (fork32_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant298_outs),
    .outs_valid (constant298_outs_valid),
    .outs_ready (constant298_outs_ready)
  );

  source source11(
    .clk (clk),
    .rst (rst),
    .outs_valid (source11_outs_valid),
    .outs_ready (source11_outs_ready)
  );

  handshake_constant_77 #(.DATA_WIDTH(5)) constant492(
    .ctrl_valid (source11_outs_valid),
    .ctrl_ready (source11_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant492_outs),
    .outs_valid (constant492_outs_valid),
    .outs_ready (constant492_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi10(
    .lhs (fork31_outs_0),
    .lhs_valid (fork31_outs_0_valid),
    .lhs_ready (fork31_outs_0_ready),
    .rhs (constant492_outs),
    .rhs_valid (constant492_outs_valid),
    .rhs_ready (constant492_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi10_result),
    .result_valid (cmpi10_result_valid),
    .result_ready (cmpi10_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork33(
    .ins (cmpi10_result),
    .ins_valid (cmpi10_result_valid),
    .ins_ready (cmpi10_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork33_outs_8, fork33_outs_7, fork33_outs_6, fork33_outs_5, fork33_outs_4, fork33_outs_3, fork33_outs_2, fork33_outs_1, fork33_outs_0}),
    .outs_valid ({fork33_outs_8_valid, fork33_outs_7_valid, fork33_outs_6_valid, fork33_outs_5_valid, fork33_outs_4_valid, fork33_outs_3_valid, fork33_outs_2_valid, fork33_outs_1_valid, fork33_outs_0_valid}),
    .outs_ready ({fork33_outs_8_ready, fork33_outs_7_ready, fork33_outs_6_ready, fork33_outs_5_ready, fork33_outs_4_ready, fork33_outs_3_ready, fork33_outs_2_ready, fork33_outs_1_ready, fork33_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br122(
    .condition (fork33_outs_4),
    .condition_valid (fork33_outs_4_valid),
    .condition_ready (fork33_outs_4_ready),
    .data (constant293_outs),
    .data_valid (constant293_outs_valid),
    .data_ready (constant293_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br122_trueOut),
    .trueOut_valid (cond_br122_trueOut_valid),
    .trueOut_ready (cond_br122_trueOut_ready),
    .falseOut (cond_br122_falseOut),
    .falseOut_valid (cond_br122_falseOut_valid),
    .falseOut_ready (cond_br122_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink80(
    .ins (cond_br122_falseOut),
    .ins_valid (cond_br122_falseOut_valid),
    .ins_ready (cond_br122_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(32)) cond_br123(
    .condition (fork33_outs_7),
    .condition_valid (fork33_outs_7_valid),
    .condition_ready (fork33_outs_7_ready),
    .data (constant489_outs),
    .data_valid (constant489_outs_valid),
    .data_ready (constant489_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br123_trueOut),
    .trueOut_valid (cond_br123_trueOut_valid),
    .trueOut_ready (cond_br123_trueOut_ready),
    .falseOut (cond_br123_falseOut),
    .falseOut_valid (cond_br123_falseOut_valid),
    .falseOut_ready (cond_br123_falseOut_ready)
  );

  sink #(.DATA_TYPE(32)) sink81(
    .ins (cond_br123_falseOut),
    .ins_valid (cond_br123_falseOut_valid),
    .ins_ready (cond_br123_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(32), .OUTPUT_TYPE(33)) extsi168(
    .ins (cond_br123_trueOut),
    .ins_valid (cond_br123_trueOut_valid),
    .ins_ready (cond_br123_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi168_outs),
    .outs_valid (extsi168_outs_valid),
    .outs_ready (extsi168_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br124(
    .condition (fork33_outs_3),
    .condition_valid (fork33_outs_3_valid),
    .condition_ready (fork33_outs_3_ready),
    .data (constant295_outs),
    .data_valid (constant295_outs_valid),
    .data_ready (constant295_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br124_trueOut),
    .trueOut_valid (cond_br124_trueOut_valid),
    .trueOut_ready (cond_br124_trueOut_ready),
    .falseOut (cond_br124_falseOut),
    .falseOut_valid (cond_br124_falseOut_valid),
    .falseOut_ready (cond_br124_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink82(
    .ins (cond_br124_falseOut),
    .ins_valid (cond_br124_falseOut_valid),
    .ins_ready (cond_br124_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(21)) cond_br125(
    .condition (fork33_outs_6),
    .condition_valid (fork33_outs_6_valid),
    .condition_ready (fork33_outs_6_ready),
    .data (constant490_outs),
    .data_valid (constant490_outs_valid),
    .data_ready (constant490_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br125_trueOut),
    .trueOut_valid (cond_br125_trueOut_valid),
    .trueOut_ready (cond_br125_trueOut_ready),
    .falseOut (cond_br125_falseOut),
    .falseOut_valid (cond_br125_falseOut_valid),
    .falseOut_ready (cond_br125_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink83(
    .ins (cond_br125_falseOut),
    .ins_valid (cond_br125_falseOut_valid),
    .ins_ready (cond_br125_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(21), .OUTPUT_TYPE(22)) extsi169(
    .ins (cond_br125_trueOut),
    .ins_valid (cond_br125_trueOut_valid),
    .ins_ready (cond_br125_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi169_outs),
    .outs_valid (extsi169_outs_valid),
    .outs_ready (extsi169_outs_ready)
  );

  cond_br #(.DATA_TYPE(15)) cond_br126(
    .condition (fork33_outs_5),
    .condition_valid (fork33_outs_5_valid),
    .condition_ready (fork33_outs_5_ready),
    .data (constant491_outs),
    .data_valid (constant491_outs_valid),
    .data_ready (constant491_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br126_trueOut),
    .trueOut_valid (cond_br126_trueOut_valid),
    .trueOut_ready (cond_br126_trueOut_ready),
    .falseOut (cond_br126_falseOut),
    .falseOut_valid (cond_br126_falseOut_valid),
    .falseOut_ready (cond_br126_falseOut_ready)
  );

  sink #(.DATA_TYPE(15)) sink84(
    .ins (cond_br126_falseOut),
    .ins_valid (cond_br126_falseOut_valid),
    .ins_ready (cond_br126_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(15), .OUTPUT_TYPE(17)) extsi170(
    .ins (cond_br126_trueOut),
    .ins_valid (cond_br126_trueOut_valid),
    .ins_ready (cond_br126_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi170_outs),
    .outs_valid (extsi170_outs_valid),
    .outs_ready (extsi170_outs_ready)
  );

  cond_br #(.DATA_TYPE(12)) cond_br127(
    .condition (fork33_outs_2),
    .condition_valid (fork33_outs_2_valid),
    .condition_ready (fork33_outs_2_ready),
    .data (constant298_outs),
    .data_valid (constant298_outs_valid),
    .data_ready (constant298_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br127_trueOut),
    .trueOut_valid (cond_br127_trueOut_valid),
    .trueOut_ready (cond_br127_trueOut_ready),
    .falseOut (cond_br127_falseOut),
    .falseOut_valid (cond_br127_falseOut_valid),
    .falseOut_ready (cond_br127_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink85(
    .ins (cond_br127_falseOut),
    .ins_valid (cond_br127_falseOut_valid),
    .ins_ready (cond_br127_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer54(
    .ins (cond_br119_falseOut),
    .ins_valid (cond_br119_falseOut_valid),
    .ins_ready (cond_br119_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer54_outs),
    .outs_valid (buffer54_outs_valid),
    .outs_ready (buffer54_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer55(
    .ins (buffer54_outs),
    .ins_valid (buffer54_outs_valid),
    .ins_ready (buffer54_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer55_outs),
    .outs_valid (buffer55_outs_valid),
    .outs_ready (buffer55_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br128(
    .condition (fork33_outs_0),
    .condition_valid (fork33_outs_0_valid),
    .condition_ready (fork33_outs_0_ready),
    .data (buffer55_outs),
    .data_valid (buffer55_outs_valid),
    .data_ready (buffer55_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br128_trueOut),
    .trueOut_valid (cond_br128_trueOut_valid),
    .trueOut_ready (cond_br128_trueOut_ready),
    .falseOut (cond_br128_falseOut),
    .falseOut_valid (cond_br128_falseOut_valid),
    .falseOut_ready (cond_br128_falseOut_ready)
  );

  cond_br_dataless cond_br129(
    .condition (fork33_outs_1),
    .condition_valid (fork33_outs_1_valid),
    .condition_ready (fork33_outs_1_ready),
    .data_valid (fork32_outs_6_valid),
    .data_ready (fork32_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br129_trueOut_valid),
    .trueOut_ready (cond_br129_trueOut_ready),
    .falseOut_valid (cond_br129_falseOut_valid),
    .falseOut_ready (cond_br129_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br130(
    .condition (fork33_outs_8),
    .condition_valid (fork33_outs_8_valid),
    .condition_ready (fork33_outs_8_ready),
    .data (fork31_outs_1),
    .data_valid (fork31_outs_1_valid),
    .data_ready (fork31_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br130_trueOut),
    .trueOut_valid (cond_br130_trueOut_valid),
    .trueOut_ready (cond_br130_trueOut_ready),
    .falseOut (cond_br130_falseOut),
    .falseOut_valid (cond_br130_falseOut_valid),
    .falseOut_ready (cond_br130_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink86(
    .ins (cond_br130_trueOut),
    .ins_valid (cond_br130_trueOut_valid),
    .ins_ready (cond_br130_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer62(
    .ins (cond_br130_falseOut),
    .ins_valid (cond_br130_falseOut_valid),
    .ins_ready (cond_br130_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer62_outs),
    .outs_valid (buffer62_outs_valid),
    .outs_ready (buffer62_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer63(
    .ins (buffer62_outs),
    .ins_valid (buffer62_outs_valid),
    .ins_ready (buffer62_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer63_outs),
    .outs_valid (buffer63_outs_valid),
    .outs_ready (buffer63_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork34(
    .ins (buffer63_outs),
    .ins_valid (buffer63_outs_valid),
    .ins_ready (buffer63_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork34_outs_1, fork34_outs_0}),
    .outs_valid ({fork34_outs_1_valid, fork34_outs_0_valid}),
    .outs_ready ({fork34_outs_1_ready, fork34_outs_0_ready})
  );

  oehb_dataless buffer64(
    .ins_valid (cond_br129_falseOut_valid),
    .ins_ready (cond_br129_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer64_outs_valid),
    .outs_ready (buffer64_outs_ready)
  );

  tehb_dataless buffer65(
    .ins_valid (buffer64_outs_valid),
    .ins_ready (buffer64_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer65_outs_valid),
    .outs_ready (buffer65_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork35(
    .ins_valid (buffer65_outs_valid),
    .ins_ready (buffer65_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork35_outs_6_valid, fork35_outs_5_valid, fork35_outs_4_valid, fork35_outs_3_valid, fork35_outs_2_valid, fork35_outs_1_valid, fork35_outs_0_valid}),
    .outs_ready ({fork35_outs_6_ready, fork35_outs_5_ready, fork35_outs_4_ready, fork35_outs_3_ready, fork35_outs_2_ready, fork35_outs_1_ready, fork35_outs_0_ready})
  );

  handshake_constant_78 #(.DATA_WIDTH(37)) constant300(
    .ctrl_valid (fork35_outs_5_valid),
    .ctrl_ready (fork35_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant300_outs),
    .outs_valid (constant300_outs_valid),
    .outs_ready (constant300_outs_ready)
  );

  handshake_constant_79 #(.DATA_WIDTH(31)) constant493(
    .ctrl_valid (fork35_outs_2_valid),
    .ctrl_ready (fork35_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant493_outs),
    .outs_valid (constant493_outs_valid),
    .outs_ready (constant493_outs_ready)
  );

  handshake_constant_80 #(.DATA_WIDTH(27)) constant302(
    .ctrl_valid (fork35_outs_4_valid),
    .ctrl_ready (fork35_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant302_outs),
    .outs_valid (constant302_outs_valid),
    .outs_ready (constant302_outs_ready)
  );

  handshake_constant_81 #(.DATA_WIDTH(21)) constant494(
    .ctrl_valid (fork35_outs_1_valid),
    .ctrl_ready (fork35_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant494_outs),
    .outs_valid (constant494_outs_valid),
    .outs_ready (constant494_outs_ready)
  );

  handshake_constant_82 #(.DATA_WIDTH(13)) constant495(
    .ctrl_valid (fork35_outs_0_valid),
    .ctrl_ready (fork35_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant495_outs),
    .outs_valid (constant495_outs_valid),
    .outs_ready (constant495_outs_ready)
  );

  handshake_constant_83 #(.DATA_WIDTH(12)) constant305(
    .ctrl_valid (fork35_outs_3_valid),
    .ctrl_ready (fork35_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant305_outs),
    .outs_valid (constant305_outs_valid),
    .outs_ready (constant305_outs_ready)
  );

  source source12(
    .clk (clk),
    .rst (rst),
    .outs_valid (source12_outs_valid),
    .outs_ready (source12_outs_ready)
  );

  handshake_constant_84 #(.DATA_WIDTH(5)) constant496(
    .ctrl_valid (source12_outs_valid),
    .ctrl_ready (source12_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant496_outs),
    .outs_valid (constant496_outs_valid),
    .outs_ready (constant496_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi11(
    .lhs (fork34_outs_0),
    .lhs_valid (fork34_outs_0_valid),
    .lhs_ready (fork34_outs_0_ready),
    .rhs (constant496_outs),
    .rhs_valid (constant496_outs_valid),
    .rhs_ready (constant496_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi11_result),
    .result_valid (cmpi11_result_valid),
    .result_ready (cmpi11_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork36(
    .ins (cmpi11_result),
    .ins_valid (cmpi11_result_valid),
    .ins_ready (cmpi11_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork36_outs_8, fork36_outs_7, fork36_outs_6, fork36_outs_5, fork36_outs_4, fork36_outs_3, fork36_outs_2, fork36_outs_1, fork36_outs_0}),
    .outs_valid ({fork36_outs_8_valid, fork36_outs_7_valid, fork36_outs_6_valid, fork36_outs_5_valid, fork36_outs_4_valid, fork36_outs_3_valid, fork36_outs_2_valid, fork36_outs_1_valid, fork36_outs_0_valid}),
    .outs_ready ({fork36_outs_8_ready, fork36_outs_7_ready, fork36_outs_6_ready, fork36_outs_5_ready, fork36_outs_4_ready, fork36_outs_3_ready, fork36_outs_2_ready, fork36_outs_1_ready, fork36_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br131(
    .condition (fork36_outs_4),
    .condition_valid (fork36_outs_4_valid),
    .condition_ready (fork36_outs_4_ready),
    .data (constant300_outs),
    .data_valid (constant300_outs_valid),
    .data_ready (constant300_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br131_trueOut),
    .trueOut_valid (cond_br131_trueOut_valid),
    .trueOut_ready (cond_br131_trueOut_ready),
    .falseOut (cond_br131_falseOut),
    .falseOut_valid (cond_br131_falseOut_valid),
    .falseOut_ready (cond_br131_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink88(
    .ins (cond_br131_falseOut),
    .ins_valid (cond_br131_falseOut_valid),
    .ins_ready (cond_br131_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(31)) cond_br132(
    .condition (fork36_outs_7),
    .condition_valid (fork36_outs_7_valid),
    .condition_ready (fork36_outs_7_ready),
    .data (constant493_outs),
    .data_valid (constant493_outs_valid),
    .data_ready (constant493_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br132_trueOut),
    .trueOut_valid (cond_br132_trueOut_valid),
    .trueOut_ready (cond_br132_trueOut_ready),
    .falseOut (cond_br132_falseOut),
    .falseOut_valid (cond_br132_falseOut_valid),
    .falseOut_ready (cond_br132_falseOut_ready)
  );

  sink #(.DATA_TYPE(31)) sink89(
    .ins (cond_br132_falseOut),
    .ins_valid (cond_br132_falseOut_valid),
    .ins_ready (cond_br132_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(31), .OUTPUT_TYPE(33)) extsi171(
    .ins (cond_br132_trueOut),
    .ins_valid (cond_br132_trueOut_valid),
    .ins_ready (cond_br132_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi171_outs),
    .outs_valid (extsi171_outs_valid),
    .outs_ready (extsi171_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br133(
    .condition (fork36_outs_3),
    .condition_valid (fork36_outs_3_valid),
    .condition_ready (fork36_outs_3_ready),
    .data (constant302_outs),
    .data_valid (constant302_outs_valid),
    .data_ready (constant302_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br133_trueOut),
    .trueOut_valid (cond_br133_trueOut_valid),
    .trueOut_ready (cond_br133_trueOut_ready),
    .falseOut (cond_br133_falseOut),
    .falseOut_valid (cond_br133_falseOut_valid),
    .falseOut_ready (cond_br133_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink90(
    .ins (cond_br133_falseOut),
    .ins_valid (cond_br133_falseOut_valid),
    .ins_ready (cond_br133_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(21)) cond_br134(
    .condition (fork36_outs_6),
    .condition_valid (fork36_outs_6_valid),
    .condition_ready (fork36_outs_6_ready),
    .data (constant494_outs),
    .data_valid (constant494_outs_valid),
    .data_ready (constant494_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br134_trueOut),
    .trueOut_valid (cond_br134_trueOut_valid),
    .trueOut_ready (cond_br134_trueOut_ready),
    .falseOut (cond_br134_falseOut),
    .falseOut_valid (cond_br134_falseOut_valid),
    .falseOut_ready (cond_br134_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink91(
    .ins (cond_br134_falseOut),
    .ins_valid (cond_br134_falseOut_valid),
    .ins_ready (cond_br134_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(21), .OUTPUT_TYPE(22)) extsi172(
    .ins (cond_br134_trueOut),
    .ins_valid (cond_br134_trueOut_valid),
    .ins_ready (cond_br134_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi172_outs),
    .outs_valid (extsi172_outs_valid),
    .outs_ready (extsi172_outs_ready)
  );

  cond_br #(.DATA_TYPE(13)) cond_br135(
    .condition (fork36_outs_5),
    .condition_valid (fork36_outs_5_valid),
    .condition_ready (fork36_outs_5_ready),
    .data (constant495_outs),
    .data_valid (constant495_outs_valid),
    .data_ready (constant495_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br135_trueOut),
    .trueOut_valid (cond_br135_trueOut_valid),
    .trueOut_ready (cond_br135_trueOut_ready),
    .falseOut (cond_br135_falseOut),
    .falseOut_valid (cond_br135_falseOut_valid),
    .falseOut_ready (cond_br135_falseOut_ready)
  );

  sink #(.DATA_TYPE(13)) sink92(
    .ins (cond_br135_falseOut),
    .ins_valid (cond_br135_falseOut_valid),
    .ins_ready (cond_br135_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(13), .OUTPUT_TYPE(17)) extsi173(
    .ins (cond_br135_trueOut),
    .ins_valid (cond_br135_trueOut_valid),
    .ins_ready (cond_br135_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi173_outs),
    .outs_valid (extsi173_outs_valid),
    .outs_ready (extsi173_outs_ready)
  );

  cond_br #(.DATA_TYPE(12)) cond_br136(
    .condition (fork36_outs_2),
    .condition_valid (fork36_outs_2_valid),
    .condition_ready (fork36_outs_2_ready),
    .data (constant305_outs),
    .data_valid (constant305_outs_valid),
    .data_ready (constant305_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br136_trueOut),
    .trueOut_valid (cond_br136_trueOut_valid),
    .trueOut_ready (cond_br136_trueOut_ready),
    .falseOut (cond_br136_falseOut),
    .falseOut_valid (cond_br136_falseOut_valid),
    .falseOut_ready (cond_br136_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink93(
    .ins (cond_br136_falseOut),
    .ins_valid (cond_br136_falseOut_valid),
    .ins_ready (cond_br136_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer60(
    .ins (cond_br128_falseOut),
    .ins_valid (cond_br128_falseOut_valid),
    .ins_ready (cond_br128_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer60_outs),
    .outs_valid (buffer60_outs_valid),
    .outs_ready (buffer60_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer61(
    .ins (buffer60_outs),
    .ins_valid (buffer60_outs_valid),
    .ins_ready (buffer60_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer61_outs),
    .outs_valid (buffer61_outs_valid),
    .outs_ready (buffer61_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br137(
    .condition (fork36_outs_0),
    .condition_valid (fork36_outs_0_valid),
    .condition_ready (fork36_outs_0_ready),
    .data (buffer61_outs),
    .data_valid (buffer61_outs_valid),
    .data_ready (buffer61_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br137_trueOut),
    .trueOut_valid (cond_br137_trueOut_valid),
    .trueOut_ready (cond_br137_trueOut_ready),
    .falseOut (cond_br137_falseOut),
    .falseOut_valid (cond_br137_falseOut_valid),
    .falseOut_ready (cond_br137_falseOut_ready)
  );

  cond_br_dataless cond_br138(
    .condition (fork36_outs_1),
    .condition_valid (fork36_outs_1_valid),
    .condition_ready (fork36_outs_1_ready),
    .data_valid (fork35_outs_6_valid),
    .data_ready (fork35_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br138_trueOut_valid),
    .trueOut_ready (cond_br138_trueOut_ready),
    .falseOut_valid (cond_br138_falseOut_valid),
    .falseOut_ready (cond_br138_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br139(
    .condition (fork36_outs_8),
    .condition_valid (fork36_outs_8_valid),
    .condition_ready (fork36_outs_8_ready),
    .data (fork34_outs_1),
    .data_valid (fork34_outs_1_valid),
    .data_ready (fork34_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br139_trueOut),
    .trueOut_valid (cond_br139_trueOut_valid),
    .trueOut_ready (cond_br139_trueOut_ready),
    .falseOut (cond_br139_falseOut),
    .falseOut_valid (cond_br139_falseOut_valid),
    .falseOut_ready (cond_br139_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink94(
    .ins (cond_br139_trueOut),
    .ins_valid (cond_br139_trueOut_valid),
    .ins_ready (cond_br139_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer68(
    .ins (cond_br139_falseOut),
    .ins_valid (cond_br139_falseOut_valid),
    .ins_ready (cond_br139_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer68_outs),
    .outs_valid (buffer68_outs_valid),
    .outs_ready (buffer68_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer69(
    .ins (buffer68_outs),
    .ins_valid (buffer68_outs_valid),
    .ins_ready (buffer68_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer69_outs),
    .outs_valid (buffer69_outs_valid),
    .outs_ready (buffer69_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork37(
    .ins (buffer69_outs),
    .ins_valid (buffer69_outs_valid),
    .ins_ready (buffer69_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork37_outs_1, fork37_outs_0}),
    .outs_valid ({fork37_outs_1_valid, fork37_outs_0_valid}),
    .outs_ready ({fork37_outs_1_ready, fork37_outs_0_ready})
  );

  oehb_dataless buffer70(
    .ins_valid (cond_br138_falseOut_valid),
    .ins_ready (cond_br138_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer70_outs_valid),
    .outs_ready (buffer70_outs_ready)
  );

  tehb_dataless buffer71(
    .ins_valid (buffer70_outs_valid),
    .ins_ready (buffer70_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer71_outs_valid),
    .outs_ready (buffer71_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork38(
    .ins_valid (buffer71_outs_valid),
    .ins_ready (buffer71_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork38_outs_6_valid, fork38_outs_5_valid, fork38_outs_4_valid, fork38_outs_3_valid, fork38_outs_2_valid, fork38_outs_1_valid, fork38_outs_0_valid}),
    .outs_ready ({fork38_outs_6_ready, fork38_outs_5_ready, fork38_outs_4_ready, fork38_outs_3_ready, fork38_outs_2_ready, fork38_outs_1_ready, fork38_outs_0_ready})
  );

  handshake_constant_85 #(.DATA_WIDTH(37)) constant307(
    .ctrl_valid (fork38_outs_5_valid),
    .ctrl_ready (fork38_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant307_outs),
    .outs_valid (constant307_outs_valid),
    .outs_ready (constant307_outs_ready)
  );

  handshake_constant_86 #(.DATA_WIDTH(31)) constant497(
    .ctrl_valid (fork38_outs_1_valid),
    .ctrl_ready (fork38_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant497_outs),
    .outs_valid (constant497_outs_valid),
    .outs_ready (constant497_outs_ready)
  );

  handshake_constant_87 #(.DATA_WIDTH(27)) constant309(
    .ctrl_valid (fork38_outs_4_valid),
    .ctrl_ready (fork38_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant309_outs),
    .outs_valid (constant309_outs_valid),
    .outs_ready (constant309_outs_ready)
  );

  handshake_constant_88 #(.DATA_WIDTH(21)) constant498(
    .ctrl_valid (fork38_outs_0_valid),
    .ctrl_ready (fork38_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant498_outs),
    .outs_valid (constant498_outs_valid),
    .outs_ready (constant498_outs_ready)
  );

  handshake_constant_89 #(.DATA_WIDTH(17)) constant311(
    .ctrl_valid (fork38_outs_3_valid),
    .ctrl_ready (fork38_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant311_outs),
    .outs_valid (constant311_outs_valid),
    .outs_ready (constant311_outs_ready)
  );

  handshake_constant_90 #(.DATA_WIDTH(12)) constant312(
    .ctrl_valid (fork38_outs_2_valid),
    .ctrl_ready (fork38_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant312_outs),
    .outs_valid (constant312_outs_valid),
    .outs_ready (constant312_outs_ready)
  );

  source source13(
    .clk (clk),
    .rst (rst),
    .outs_valid (source13_outs_valid),
    .outs_ready (source13_outs_ready)
  );

  handshake_constant_7 #(.DATA_WIDTH(5)) constant499(
    .ctrl_valid (source13_outs_valid),
    .ctrl_ready (source13_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant499_outs),
    .outs_valid (constant499_outs_valid),
    .outs_ready (constant499_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi12(
    .lhs (fork37_outs_0),
    .lhs_valid (fork37_outs_0_valid),
    .lhs_ready (fork37_outs_0_ready),
    .rhs (constant499_outs),
    .rhs_valid (constant499_outs_valid),
    .rhs_ready (constant499_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi12_result),
    .result_valid (cmpi12_result_valid),
    .result_ready (cmpi12_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork39(
    .ins (cmpi12_result),
    .ins_valid (cmpi12_result_valid),
    .ins_ready (cmpi12_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork39_outs_8, fork39_outs_7, fork39_outs_6, fork39_outs_5, fork39_outs_4, fork39_outs_3, fork39_outs_2, fork39_outs_1, fork39_outs_0}),
    .outs_valid ({fork39_outs_8_valid, fork39_outs_7_valid, fork39_outs_6_valid, fork39_outs_5_valid, fork39_outs_4_valid, fork39_outs_3_valid, fork39_outs_2_valid, fork39_outs_1_valid, fork39_outs_0_valid}),
    .outs_ready ({fork39_outs_8_ready, fork39_outs_7_ready, fork39_outs_6_ready, fork39_outs_5_ready, fork39_outs_4_ready, fork39_outs_3_ready, fork39_outs_2_ready, fork39_outs_1_ready, fork39_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br140(
    .condition (fork39_outs_5),
    .condition_valid (fork39_outs_5_valid),
    .condition_ready (fork39_outs_5_ready),
    .data (constant307_outs),
    .data_valid (constant307_outs_valid),
    .data_ready (constant307_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br140_trueOut),
    .trueOut_valid (cond_br140_trueOut_valid),
    .trueOut_ready (cond_br140_trueOut_ready),
    .falseOut (cond_br140_falseOut),
    .falseOut_valid (cond_br140_falseOut_valid),
    .falseOut_ready (cond_br140_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink96(
    .ins (cond_br140_falseOut),
    .ins_valid (cond_br140_falseOut_valid),
    .ins_ready (cond_br140_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(31)) cond_br141(
    .condition (fork39_outs_7),
    .condition_valid (fork39_outs_7_valid),
    .condition_ready (fork39_outs_7_ready),
    .data (constant497_outs),
    .data_valid (constant497_outs_valid),
    .data_ready (constant497_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br141_trueOut),
    .trueOut_valid (cond_br141_trueOut_valid),
    .trueOut_ready (cond_br141_trueOut_ready),
    .falseOut (cond_br141_falseOut),
    .falseOut_valid (cond_br141_falseOut_valid),
    .falseOut_ready (cond_br141_falseOut_ready)
  );

  sink #(.DATA_TYPE(31)) sink97(
    .ins (cond_br141_falseOut),
    .ins_valid (cond_br141_falseOut_valid),
    .ins_ready (cond_br141_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(31), .OUTPUT_TYPE(33)) extsi174(
    .ins (cond_br141_trueOut),
    .ins_valid (cond_br141_trueOut_valid),
    .ins_ready (cond_br141_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi174_outs),
    .outs_valid (extsi174_outs_valid),
    .outs_ready (extsi174_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br142(
    .condition (fork39_outs_4),
    .condition_valid (fork39_outs_4_valid),
    .condition_ready (fork39_outs_4_ready),
    .data (constant309_outs),
    .data_valid (constant309_outs_valid),
    .data_ready (constant309_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br142_trueOut),
    .trueOut_valid (cond_br142_trueOut_valid),
    .trueOut_ready (cond_br142_trueOut_ready),
    .falseOut (cond_br142_falseOut),
    .falseOut_valid (cond_br142_falseOut_valid),
    .falseOut_ready (cond_br142_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink98(
    .ins (cond_br142_falseOut),
    .ins_valid (cond_br142_falseOut_valid),
    .ins_ready (cond_br142_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(21)) cond_br143(
    .condition (fork39_outs_6),
    .condition_valid (fork39_outs_6_valid),
    .condition_ready (fork39_outs_6_ready),
    .data (constant498_outs),
    .data_valid (constant498_outs_valid),
    .data_ready (constant498_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br143_trueOut),
    .trueOut_valid (cond_br143_trueOut_valid),
    .trueOut_ready (cond_br143_trueOut_ready),
    .falseOut (cond_br143_falseOut),
    .falseOut_valid (cond_br143_falseOut_valid),
    .falseOut_ready (cond_br143_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink99(
    .ins (cond_br143_falseOut),
    .ins_valid (cond_br143_falseOut_valid),
    .ins_ready (cond_br143_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(21), .OUTPUT_TYPE(22)) extsi175(
    .ins (cond_br143_trueOut),
    .ins_valid (cond_br143_trueOut_valid),
    .ins_ready (cond_br143_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi175_outs),
    .outs_valid (extsi175_outs_valid),
    .outs_ready (extsi175_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br144(
    .condition (fork39_outs_3),
    .condition_valid (fork39_outs_3_valid),
    .condition_ready (fork39_outs_3_ready),
    .data (constant311_outs),
    .data_valid (constant311_outs_valid),
    .data_ready (constant311_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br144_trueOut),
    .trueOut_valid (cond_br144_trueOut_valid),
    .trueOut_ready (cond_br144_trueOut_ready),
    .falseOut (cond_br144_falseOut),
    .falseOut_valid (cond_br144_falseOut_valid),
    .falseOut_ready (cond_br144_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink100(
    .ins (cond_br144_falseOut),
    .ins_valid (cond_br144_falseOut_valid),
    .ins_ready (cond_br144_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br145(
    .condition (fork39_outs_2),
    .condition_valid (fork39_outs_2_valid),
    .condition_ready (fork39_outs_2_ready),
    .data (constant312_outs),
    .data_valid (constant312_outs_valid),
    .data_ready (constant312_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br145_trueOut),
    .trueOut_valid (cond_br145_trueOut_valid),
    .trueOut_ready (cond_br145_trueOut_ready),
    .falseOut (cond_br145_falseOut),
    .falseOut_valid (cond_br145_falseOut_valid),
    .falseOut_ready (cond_br145_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink101(
    .ins (cond_br145_falseOut),
    .ins_valid (cond_br145_falseOut_valid),
    .ins_ready (cond_br145_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer66(
    .ins (cond_br137_falseOut),
    .ins_valid (cond_br137_falseOut_valid),
    .ins_ready (cond_br137_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer66_outs),
    .outs_valid (buffer66_outs_valid),
    .outs_ready (buffer66_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer67(
    .ins (buffer66_outs),
    .ins_valid (buffer66_outs_valid),
    .ins_ready (buffer66_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer67_outs),
    .outs_valid (buffer67_outs_valid),
    .outs_ready (buffer67_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br146(
    .condition (fork39_outs_0),
    .condition_valid (fork39_outs_0_valid),
    .condition_ready (fork39_outs_0_ready),
    .data (buffer67_outs),
    .data_valid (buffer67_outs_valid),
    .data_ready (buffer67_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br146_trueOut),
    .trueOut_valid (cond_br146_trueOut_valid),
    .trueOut_ready (cond_br146_trueOut_ready),
    .falseOut (cond_br146_falseOut),
    .falseOut_valid (cond_br146_falseOut_valid),
    .falseOut_ready (cond_br146_falseOut_ready)
  );

  cond_br_dataless cond_br147(
    .condition (fork39_outs_1),
    .condition_valid (fork39_outs_1_valid),
    .condition_ready (fork39_outs_1_ready),
    .data_valid (fork38_outs_6_valid),
    .data_ready (fork38_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br147_trueOut_valid),
    .trueOut_ready (cond_br147_trueOut_ready),
    .falseOut_valid (cond_br147_falseOut_valid),
    .falseOut_ready (cond_br147_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br148(
    .condition (fork39_outs_8),
    .condition_valid (fork39_outs_8_valid),
    .condition_ready (fork39_outs_8_ready),
    .data (fork37_outs_1),
    .data_valid (fork37_outs_1_valid),
    .data_ready (fork37_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br148_trueOut),
    .trueOut_valid (cond_br148_trueOut_valid),
    .trueOut_ready (cond_br148_trueOut_ready),
    .falseOut (cond_br148_falseOut),
    .falseOut_valid (cond_br148_falseOut_valid),
    .falseOut_ready (cond_br148_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink102(
    .ins (cond_br148_trueOut),
    .ins_valid (cond_br148_trueOut_valid),
    .ins_ready (cond_br148_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer74(
    .ins (cond_br148_falseOut),
    .ins_valid (cond_br148_falseOut_valid),
    .ins_ready (cond_br148_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer74_outs),
    .outs_valid (buffer74_outs_valid),
    .outs_ready (buffer74_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer75(
    .ins (buffer74_outs),
    .ins_valid (buffer74_outs_valid),
    .ins_ready (buffer74_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer75_outs),
    .outs_valid (buffer75_outs_valid),
    .outs_ready (buffer75_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork40(
    .ins (buffer75_outs),
    .ins_valid (buffer75_outs_valid),
    .ins_ready (buffer75_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork40_outs_1, fork40_outs_0}),
    .outs_valid ({fork40_outs_1_valid, fork40_outs_0_valid}),
    .outs_ready ({fork40_outs_1_ready, fork40_outs_0_ready})
  );

  oehb_dataless buffer76(
    .ins_valid (cond_br147_falseOut_valid),
    .ins_ready (cond_br147_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer76_outs_valid),
    .outs_ready (buffer76_outs_ready)
  );

  tehb_dataless buffer77(
    .ins_valid (buffer76_outs_valid),
    .ins_ready (buffer76_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer77_outs_valid),
    .outs_ready (buffer77_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork41(
    .ins_valid (buffer77_outs_valid),
    .ins_ready (buffer77_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork41_outs_6_valid, fork41_outs_5_valid, fork41_outs_4_valid, fork41_outs_3_valid, fork41_outs_2_valid, fork41_outs_1_valid, fork41_outs_0_valid}),
    .outs_ready ({fork41_outs_6_ready, fork41_outs_5_ready, fork41_outs_4_ready, fork41_outs_3_ready, fork41_outs_2_ready, fork41_outs_1_ready, fork41_outs_0_ready})
  );

  handshake_constant_91 #(.DATA_WIDTH(37)) constant314(
    .ctrl_valid (fork41_outs_5_valid),
    .ctrl_ready (fork41_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant314_outs),
    .outs_valid (constant314_outs_valid),
    .outs_ready (constant314_outs_ready)
  );

  handshake_constant_92 #(.DATA_WIDTH(31)) constant500(
    .ctrl_valid (fork41_outs_1_valid),
    .ctrl_ready (fork41_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant500_outs),
    .outs_valid (constant500_outs_valid),
    .outs_ready (constant500_outs_ready)
  );

  handshake_constant_93 #(.DATA_WIDTH(27)) constant316(
    .ctrl_valid (fork41_outs_4_valid),
    .ctrl_ready (fork41_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant316_outs),
    .outs_valid (constant316_outs_valid),
    .outs_ready (constant316_outs_ready)
  );

  handshake_constant_94 #(.DATA_WIDTH(21)) constant501(
    .ctrl_valid (fork41_outs_0_valid),
    .ctrl_ready (fork41_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant501_outs),
    .outs_valid (constant501_outs_valid),
    .outs_ready (constant501_outs_ready)
  );

  handshake_constant_95 #(.DATA_WIDTH(17)) constant318(
    .ctrl_valid (fork41_outs_3_valid),
    .ctrl_ready (fork41_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant318_outs),
    .outs_valid (constant318_outs_valid),
    .outs_ready (constant318_outs_ready)
  );

  handshake_constant_96 #(.DATA_WIDTH(12)) constant319(
    .ctrl_valid (fork41_outs_2_valid),
    .ctrl_ready (fork41_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant319_outs),
    .outs_valid (constant319_outs_valid),
    .outs_ready (constant319_outs_ready)
  );

  source source14(
    .clk (clk),
    .rst (rst),
    .outs_valid (source14_outs_valid),
    .outs_ready (source14_outs_ready)
  );

  handshake_constant_97 #(.DATA_WIDTH(5)) constant502(
    .ctrl_valid (source14_outs_valid),
    .ctrl_ready (source14_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant502_outs),
    .outs_valid (constant502_outs_valid),
    .outs_ready (constant502_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi13(
    .lhs (fork40_outs_0),
    .lhs_valid (fork40_outs_0_valid),
    .lhs_ready (fork40_outs_0_ready),
    .rhs (constant502_outs),
    .rhs_valid (constant502_outs_valid),
    .rhs_ready (constant502_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi13_result),
    .result_valid (cmpi13_result_valid),
    .result_ready (cmpi13_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork42(
    .ins (cmpi13_result),
    .ins_valid (cmpi13_result_valid),
    .ins_ready (cmpi13_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork42_outs_8, fork42_outs_7, fork42_outs_6, fork42_outs_5, fork42_outs_4, fork42_outs_3, fork42_outs_2, fork42_outs_1, fork42_outs_0}),
    .outs_valid ({fork42_outs_8_valid, fork42_outs_7_valid, fork42_outs_6_valid, fork42_outs_5_valid, fork42_outs_4_valid, fork42_outs_3_valid, fork42_outs_2_valid, fork42_outs_1_valid, fork42_outs_0_valid}),
    .outs_ready ({fork42_outs_8_ready, fork42_outs_7_ready, fork42_outs_6_ready, fork42_outs_5_ready, fork42_outs_4_ready, fork42_outs_3_ready, fork42_outs_2_ready, fork42_outs_1_ready, fork42_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br149(
    .condition (fork42_outs_5),
    .condition_valid (fork42_outs_5_valid),
    .condition_ready (fork42_outs_5_ready),
    .data (constant314_outs),
    .data_valid (constant314_outs_valid),
    .data_ready (constant314_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br149_trueOut),
    .trueOut_valid (cond_br149_trueOut_valid),
    .trueOut_ready (cond_br149_trueOut_ready),
    .falseOut (cond_br149_falseOut),
    .falseOut_valid (cond_br149_falseOut_valid),
    .falseOut_ready (cond_br149_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink104(
    .ins (cond_br149_falseOut),
    .ins_valid (cond_br149_falseOut_valid),
    .ins_ready (cond_br149_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(31)) cond_br150(
    .condition (fork42_outs_7),
    .condition_valid (fork42_outs_7_valid),
    .condition_ready (fork42_outs_7_ready),
    .data (constant500_outs),
    .data_valid (constant500_outs_valid),
    .data_ready (constant500_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br150_trueOut),
    .trueOut_valid (cond_br150_trueOut_valid),
    .trueOut_ready (cond_br150_trueOut_ready),
    .falseOut (cond_br150_falseOut),
    .falseOut_valid (cond_br150_falseOut_valid),
    .falseOut_ready (cond_br150_falseOut_ready)
  );

  sink #(.DATA_TYPE(31)) sink105(
    .ins (cond_br150_falseOut),
    .ins_valid (cond_br150_falseOut_valid),
    .ins_ready (cond_br150_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(31), .OUTPUT_TYPE(33)) extsi176(
    .ins (cond_br150_trueOut),
    .ins_valid (cond_br150_trueOut_valid),
    .ins_ready (cond_br150_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi176_outs),
    .outs_valid (extsi176_outs_valid),
    .outs_ready (extsi176_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br151(
    .condition (fork42_outs_4),
    .condition_valid (fork42_outs_4_valid),
    .condition_ready (fork42_outs_4_ready),
    .data (constant316_outs),
    .data_valid (constant316_outs_valid),
    .data_ready (constant316_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br151_trueOut),
    .trueOut_valid (cond_br151_trueOut_valid),
    .trueOut_ready (cond_br151_trueOut_ready),
    .falseOut (cond_br151_falseOut),
    .falseOut_valid (cond_br151_falseOut_valid),
    .falseOut_ready (cond_br151_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink106(
    .ins (cond_br151_falseOut),
    .ins_valid (cond_br151_falseOut_valid),
    .ins_ready (cond_br151_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(21)) cond_br152(
    .condition (fork42_outs_6),
    .condition_valid (fork42_outs_6_valid),
    .condition_ready (fork42_outs_6_ready),
    .data (constant501_outs),
    .data_valid (constant501_outs_valid),
    .data_ready (constant501_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br152_trueOut),
    .trueOut_valid (cond_br152_trueOut_valid),
    .trueOut_ready (cond_br152_trueOut_ready),
    .falseOut (cond_br152_falseOut),
    .falseOut_valid (cond_br152_falseOut_valid),
    .falseOut_ready (cond_br152_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink107(
    .ins (cond_br152_falseOut),
    .ins_valid (cond_br152_falseOut_valid),
    .ins_ready (cond_br152_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(21), .OUTPUT_TYPE(22)) extsi177(
    .ins (cond_br152_trueOut),
    .ins_valid (cond_br152_trueOut_valid),
    .ins_ready (cond_br152_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi177_outs),
    .outs_valid (extsi177_outs_valid),
    .outs_ready (extsi177_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br153(
    .condition (fork42_outs_3),
    .condition_valid (fork42_outs_3_valid),
    .condition_ready (fork42_outs_3_ready),
    .data (constant318_outs),
    .data_valid (constant318_outs_valid),
    .data_ready (constant318_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br153_trueOut),
    .trueOut_valid (cond_br153_trueOut_valid),
    .trueOut_ready (cond_br153_trueOut_ready),
    .falseOut (cond_br153_falseOut),
    .falseOut_valid (cond_br153_falseOut_valid),
    .falseOut_ready (cond_br153_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink108(
    .ins (cond_br153_falseOut),
    .ins_valid (cond_br153_falseOut_valid),
    .ins_ready (cond_br153_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br154(
    .condition (fork42_outs_2),
    .condition_valid (fork42_outs_2_valid),
    .condition_ready (fork42_outs_2_ready),
    .data (constant319_outs),
    .data_valid (constant319_outs_valid),
    .data_ready (constant319_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br154_trueOut),
    .trueOut_valid (cond_br154_trueOut_valid),
    .trueOut_ready (cond_br154_trueOut_ready),
    .falseOut (cond_br154_falseOut),
    .falseOut_valid (cond_br154_falseOut_valid),
    .falseOut_ready (cond_br154_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink109(
    .ins (cond_br154_falseOut),
    .ins_valid (cond_br154_falseOut_valid),
    .ins_ready (cond_br154_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer72(
    .ins (cond_br146_falseOut),
    .ins_valid (cond_br146_falseOut_valid),
    .ins_ready (cond_br146_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer72_outs),
    .outs_valid (buffer72_outs_valid),
    .outs_ready (buffer72_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer73(
    .ins (buffer72_outs),
    .ins_valid (buffer72_outs_valid),
    .ins_ready (buffer72_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer73_outs),
    .outs_valid (buffer73_outs_valid),
    .outs_ready (buffer73_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br155(
    .condition (fork42_outs_0),
    .condition_valid (fork42_outs_0_valid),
    .condition_ready (fork42_outs_0_ready),
    .data (buffer73_outs),
    .data_valid (buffer73_outs_valid),
    .data_ready (buffer73_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br155_trueOut),
    .trueOut_valid (cond_br155_trueOut_valid),
    .trueOut_ready (cond_br155_trueOut_ready),
    .falseOut (cond_br155_falseOut),
    .falseOut_valid (cond_br155_falseOut_valid),
    .falseOut_ready (cond_br155_falseOut_ready)
  );

  cond_br_dataless cond_br156(
    .condition (fork42_outs_1),
    .condition_valid (fork42_outs_1_valid),
    .condition_ready (fork42_outs_1_ready),
    .data_valid (fork41_outs_6_valid),
    .data_ready (fork41_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br156_trueOut_valid),
    .trueOut_ready (cond_br156_trueOut_ready),
    .falseOut_valid (cond_br156_falseOut_valid),
    .falseOut_ready (cond_br156_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br157(
    .condition (fork42_outs_8),
    .condition_valid (fork42_outs_8_valid),
    .condition_ready (fork42_outs_8_ready),
    .data (fork40_outs_1),
    .data_valid (fork40_outs_1_valid),
    .data_ready (fork40_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br157_trueOut),
    .trueOut_valid (cond_br157_trueOut_valid),
    .trueOut_ready (cond_br157_trueOut_ready),
    .falseOut (cond_br157_falseOut),
    .falseOut_valid (cond_br157_falseOut_valid),
    .falseOut_ready (cond_br157_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink110(
    .ins (cond_br157_trueOut),
    .ins_valid (cond_br157_trueOut_valid),
    .ins_ready (cond_br157_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer80(
    .ins (cond_br157_falseOut),
    .ins_valid (cond_br157_falseOut_valid),
    .ins_ready (cond_br157_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer80_outs),
    .outs_valid (buffer80_outs_valid),
    .outs_ready (buffer80_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer81(
    .ins (buffer80_outs),
    .ins_valid (buffer80_outs_valid),
    .ins_ready (buffer80_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer81_outs),
    .outs_valid (buffer81_outs_valid),
    .outs_ready (buffer81_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork43(
    .ins (buffer81_outs),
    .ins_valid (buffer81_outs_valid),
    .ins_ready (buffer81_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork43_outs_1, fork43_outs_0}),
    .outs_valid ({fork43_outs_1_valid, fork43_outs_0_valid}),
    .outs_ready ({fork43_outs_1_ready, fork43_outs_0_ready})
  );

  oehb_dataless buffer82(
    .ins_valid (cond_br156_falseOut_valid),
    .ins_ready (cond_br156_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer82_outs_valid),
    .outs_ready (buffer82_outs_ready)
  );

  tehb_dataless buffer83(
    .ins_valid (buffer82_outs_valid),
    .ins_ready (buffer82_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer83_outs_valid),
    .outs_ready (buffer83_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork44(
    .ins_valid (buffer83_outs_valid),
    .ins_ready (buffer83_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork44_outs_6_valid, fork44_outs_5_valid, fork44_outs_4_valid, fork44_outs_3_valid, fork44_outs_2_valid, fork44_outs_1_valid, fork44_outs_0_valid}),
    .outs_ready ({fork44_outs_6_ready, fork44_outs_5_ready, fork44_outs_4_ready, fork44_outs_3_ready, fork44_outs_2_ready, fork44_outs_1_ready, fork44_outs_0_ready})
  );

  handshake_constant_98 #(.DATA_WIDTH(37)) constant321(
    .ctrl_valid (fork44_outs_5_valid),
    .ctrl_ready (fork44_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant321_outs),
    .outs_valid (constant321_outs_valid),
    .outs_ready (constant321_outs_ready)
  );

  handshake_constant_99 #(.DATA_WIDTH(31)) constant503(
    .ctrl_valid (fork44_outs_1_valid),
    .ctrl_ready (fork44_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant503_outs),
    .outs_valid (constant503_outs_valid),
    .outs_ready (constant503_outs_ready)
  );

  handshake_constant_100 #(.DATA_WIDTH(27)) constant323(
    .ctrl_valid (fork44_outs_4_valid),
    .ctrl_ready (fork44_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant323_outs),
    .outs_valid (constant323_outs_valid),
    .outs_ready (constant323_outs_ready)
  );

  handshake_constant_101 #(.DATA_WIDTH(21)) constant504(
    .ctrl_valid (fork44_outs_0_valid),
    .ctrl_ready (fork44_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant504_outs),
    .outs_valid (constant504_outs_valid),
    .outs_ready (constant504_outs_ready)
  );

  handshake_constant_102 #(.DATA_WIDTH(17)) constant325(
    .ctrl_valid (fork44_outs_3_valid),
    .ctrl_ready (fork44_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant325_outs),
    .outs_valid (constant325_outs_valid),
    .outs_ready (constant325_outs_ready)
  );

  handshake_constant_103 #(.DATA_WIDTH(12)) constant326(
    .ctrl_valid (fork44_outs_2_valid),
    .ctrl_ready (fork44_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant326_outs),
    .outs_valid (constant326_outs_valid),
    .outs_ready (constant326_outs_ready)
  );

  source source15(
    .clk (clk),
    .rst (rst),
    .outs_valid (source15_outs_valid),
    .outs_ready (source15_outs_ready)
  );

  handshake_constant_104 #(.DATA_WIDTH(5)) constant505(
    .ctrl_valid (source15_outs_valid),
    .ctrl_ready (source15_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant505_outs),
    .outs_valid (constant505_outs_valid),
    .outs_ready (constant505_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi14(
    .lhs (fork43_outs_0),
    .lhs_valid (fork43_outs_0_valid),
    .lhs_ready (fork43_outs_0_ready),
    .rhs (constant505_outs),
    .rhs_valid (constant505_outs_valid),
    .rhs_ready (constant505_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi14_result),
    .result_valid (cmpi14_result_valid),
    .result_ready (cmpi14_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork45(
    .ins (cmpi14_result),
    .ins_valid (cmpi14_result_valid),
    .ins_ready (cmpi14_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork45_outs_8, fork45_outs_7, fork45_outs_6, fork45_outs_5, fork45_outs_4, fork45_outs_3, fork45_outs_2, fork45_outs_1, fork45_outs_0}),
    .outs_valid ({fork45_outs_8_valid, fork45_outs_7_valid, fork45_outs_6_valid, fork45_outs_5_valid, fork45_outs_4_valid, fork45_outs_3_valid, fork45_outs_2_valid, fork45_outs_1_valid, fork45_outs_0_valid}),
    .outs_ready ({fork45_outs_8_ready, fork45_outs_7_ready, fork45_outs_6_ready, fork45_outs_5_ready, fork45_outs_4_ready, fork45_outs_3_ready, fork45_outs_2_ready, fork45_outs_1_ready, fork45_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br158(
    .condition (fork45_outs_5),
    .condition_valid (fork45_outs_5_valid),
    .condition_ready (fork45_outs_5_ready),
    .data (constant321_outs),
    .data_valid (constant321_outs_valid),
    .data_ready (constant321_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br158_trueOut),
    .trueOut_valid (cond_br158_trueOut_valid),
    .trueOut_ready (cond_br158_trueOut_ready),
    .falseOut (cond_br158_falseOut),
    .falseOut_valid (cond_br158_falseOut_valid),
    .falseOut_ready (cond_br158_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink112(
    .ins (cond_br158_falseOut),
    .ins_valid (cond_br158_falseOut_valid),
    .ins_ready (cond_br158_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(31)) cond_br159(
    .condition (fork45_outs_7),
    .condition_valid (fork45_outs_7_valid),
    .condition_ready (fork45_outs_7_ready),
    .data (constant503_outs),
    .data_valid (constant503_outs_valid),
    .data_ready (constant503_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br159_trueOut),
    .trueOut_valid (cond_br159_trueOut_valid),
    .trueOut_ready (cond_br159_trueOut_ready),
    .falseOut (cond_br159_falseOut),
    .falseOut_valid (cond_br159_falseOut_valid),
    .falseOut_ready (cond_br159_falseOut_ready)
  );

  sink #(.DATA_TYPE(31)) sink113(
    .ins (cond_br159_falseOut),
    .ins_valid (cond_br159_falseOut_valid),
    .ins_ready (cond_br159_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(31), .OUTPUT_TYPE(33)) extsi178(
    .ins (cond_br159_trueOut),
    .ins_valid (cond_br159_trueOut_valid),
    .ins_ready (cond_br159_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi178_outs),
    .outs_valid (extsi178_outs_valid),
    .outs_ready (extsi178_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br160(
    .condition (fork45_outs_4),
    .condition_valid (fork45_outs_4_valid),
    .condition_ready (fork45_outs_4_ready),
    .data (constant323_outs),
    .data_valid (constant323_outs_valid),
    .data_ready (constant323_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br160_trueOut),
    .trueOut_valid (cond_br160_trueOut_valid),
    .trueOut_ready (cond_br160_trueOut_ready),
    .falseOut (cond_br160_falseOut),
    .falseOut_valid (cond_br160_falseOut_valid),
    .falseOut_ready (cond_br160_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink114(
    .ins (cond_br160_falseOut),
    .ins_valid (cond_br160_falseOut_valid),
    .ins_ready (cond_br160_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(21)) cond_br161(
    .condition (fork45_outs_6),
    .condition_valid (fork45_outs_6_valid),
    .condition_ready (fork45_outs_6_ready),
    .data (constant504_outs),
    .data_valid (constant504_outs_valid),
    .data_ready (constant504_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br161_trueOut),
    .trueOut_valid (cond_br161_trueOut_valid),
    .trueOut_ready (cond_br161_trueOut_ready),
    .falseOut (cond_br161_falseOut),
    .falseOut_valid (cond_br161_falseOut_valid),
    .falseOut_ready (cond_br161_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink115(
    .ins (cond_br161_falseOut),
    .ins_valid (cond_br161_falseOut_valid),
    .ins_ready (cond_br161_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(21), .OUTPUT_TYPE(22)) extsi179(
    .ins (cond_br161_trueOut),
    .ins_valid (cond_br161_trueOut_valid),
    .ins_ready (cond_br161_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi179_outs),
    .outs_valid (extsi179_outs_valid),
    .outs_ready (extsi179_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br162(
    .condition (fork45_outs_3),
    .condition_valid (fork45_outs_3_valid),
    .condition_ready (fork45_outs_3_ready),
    .data (constant325_outs),
    .data_valid (constant325_outs_valid),
    .data_ready (constant325_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br162_trueOut),
    .trueOut_valid (cond_br162_trueOut_valid),
    .trueOut_ready (cond_br162_trueOut_ready),
    .falseOut (cond_br162_falseOut),
    .falseOut_valid (cond_br162_falseOut_valid),
    .falseOut_ready (cond_br162_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink116(
    .ins (cond_br162_falseOut),
    .ins_valid (cond_br162_falseOut_valid),
    .ins_ready (cond_br162_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br163(
    .condition (fork45_outs_2),
    .condition_valid (fork45_outs_2_valid),
    .condition_ready (fork45_outs_2_ready),
    .data (constant326_outs),
    .data_valid (constant326_outs_valid),
    .data_ready (constant326_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br163_trueOut),
    .trueOut_valid (cond_br163_trueOut_valid),
    .trueOut_ready (cond_br163_trueOut_ready),
    .falseOut (cond_br163_falseOut),
    .falseOut_valid (cond_br163_falseOut_valid),
    .falseOut_ready (cond_br163_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink117(
    .ins (cond_br163_falseOut),
    .ins_valid (cond_br163_falseOut_valid),
    .ins_ready (cond_br163_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer78(
    .ins (cond_br155_falseOut),
    .ins_valid (cond_br155_falseOut_valid),
    .ins_ready (cond_br155_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer78_outs),
    .outs_valid (buffer78_outs_valid),
    .outs_ready (buffer78_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer79(
    .ins (buffer78_outs),
    .ins_valid (buffer78_outs_valid),
    .ins_ready (buffer78_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer79_outs),
    .outs_valid (buffer79_outs_valid),
    .outs_ready (buffer79_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br164(
    .condition (fork45_outs_0),
    .condition_valid (fork45_outs_0_valid),
    .condition_ready (fork45_outs_0_ready),
    .data (buffer79_outs),
    .data_valid (buffer79_outs_valid),
    .data_ready (buffer79_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br164_trueOut),
    .trueOut_valid (cond_br164_trueOut_valid),
    .trueOut_ready (cond_br164_trueOut_ready),
    .falseOut (cond_br164_falseOut),
    .falseOut_valid (cond_br164_falseOut_valid),
    .falseOut_ready (cond_br164_falseOut_ready)
  );

  cond_br_dataless cond_br165(
    .condition (fork45_outs_1),
    .condition_valid (fork45_outs_1_valid),
    .condition_ready (fork45_outs_1_ready),
    .data_valid (fork44_outs_6_valid),
    .data_ready (fork44_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br165_trueOut_valid),
    .trueOut_ready (cond_br165_trueOut_ready),
    .falseOut_valid (cond_br165_falseOut_valid),
    .falseOut_ready (cond_br165_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br166(
    .condition (fork45_outs_8),
    .condition_valid (fork45_outs_8_valid),
    .condition_ready (fork45_outs_8_ready),
    .data (fork43_outs_1),
    .data_valid (fork43_outs_1_valid),
    .data_ready (fork43_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br166_trueOut),
    .trueOut_valid (cond_br166_trueOut_valid),
    .trueOut_ready (cond_br166_trueOut_ready),
    .falseOut (cond_br166_falseOut),
    .falseOut_valid (cond_br166_falseOut_valid),
    .falseOut_ready (cond_br166_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink118(
    .ins (cond_br166_trueOut),
    .ins_valid (cond_br166_trueOut_valid),
    .ins_ready (cond_br166_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer86(
    .ins (cond_br166_falseOut),
    .ins_valid (cond_br166_falseOut_valid),
    .ins_ready (cond_br166_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer86_outs),
    .outs_valid (buffer86_outs_valid),
    .outs_ready (buffer86_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer87(
    .ins (buffer86_outs),
    .ins_valid (buffer86_outs_valid),
    .ins_ready (buffer86_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer87_outs),
    .outs_valid (buffer87_outs_valid),
    .outs_ready (buffer87_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork46(
    .ins (buffer87_outs),
    .ins_valid (buffer87_outs_valid),
    .ins_ready (buffer87_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork46_outs_1, fork46_outs_0}),
    .outs_valid ({fork46_outs_1_valid, fork46_outs_0_valid}),
    .outs_ready ({fork46_outs_1_ready, fork46_outs_0_ready})
  );

  oehb_dataless buffer88(
    .ins_valid (cond_br165_falseOut_valid),
    .ins_ready (cond_br165_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer88_outs_valid),
    .outs_ready (buffer88_outs_ready)
  );

  tehb_dataless buffer89(
    .ins_valid (buffer88_outs_valid),
    .ins_ready (buffer88_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer89_outs_valid),
    .outs_ready (buffer89_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork47(
    .ins_valid (buffer89_outs_valid),
    .ins_ready (buffer89_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork47_outs_6_valid, fork47_outs_5_valid, fork47_outs_4_valid, fork47_outs_3_valid, fork47_outs_2_valid, fork47_outs_1_valid, fork47_outs_0_valid}),
    .outs_ready ({fork47_outs_6_ready, fork47_outs_5_ready, fork47_outs_4_ready, fork47_outs_3_ready, fork47_outs_2_ready, fork47_outs_1_ready, fork47_outs_0_ready})
  );

  handshake_constant_105 #(.DATA_WIDTH(37)) constant328(
    .ctrl_valid (fork47_outs_5_valid),
    .ctrl_ready (fork47_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant328_outs),
    .outs_valid (constant328_outs_valid),
    .outs_ready (constant328_outs_ready)
  );

  handshake_constant_106 #(.DATA_WIDTH(31)) constant506(
    .ctrl_valid (fork47_outs_1_valid),
    .ctrl_ready (fork47_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant506_outs),
    .outs_valid (constant506_outs_valid),
    .outs_ready (constant506_outs_ready)
  );

  handshake_constant_107 #(.DATA_WIDTH(27)) constant330(
    .ctrl_valid (fork47_outs_4_valid),
    .ctrl_ready (fork47_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant330_outs),
    .outs_valid (constant330_outs_valid),
    .outs_ready (constant330_outs_ready)
  );

  handshake_constant_108 #(.DATA_WIDTH(21)) constant507(
    .ctrl_valid (fork47_outs_0_valid),
    .ctrl_ready (fork47_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant507_outs),
    .outs_valid (constant507_outs_valid),
    .outs_ready (constant507_outs_ready)
  );

  handshake_constant_109 #(.DATA_WIDTH(17)) constant332(
    .ctrl_valid (fork47_outs_3_valid),
    .ctrl_ready (fork47_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant332_outs),
    .outs_valid (constant332_outs_valid),
    .outs_ready (constant332_outs_ready)
  );

  handshake_constant_110 #(.DATA_WIDTH(12)) constant333(
    .ctrl_valid (fork47_outs_2_valid),
    .ctrl_ready (fork47_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant333_outs),
    .outs_valid (constant333_outs_valid),
    .outs_ready (constant333_outs_ready)
  );

  source source16(
    .clk (clk),
    .rst (rst),
    .outs_valid (source16_outs_valid),
    .outs_ready (source16_outs_ready)
  );

  handshake_constant_111 #(.DATA_WIDTH(5)) constant508(
    .ctrl_valid (source16_outs_valid),
    .ctrl_ready (source16_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant508_outs),
    .outs_valid (constant508_outs_valid),
    .outs_ready (constant508_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(5)) cmpi15(
    .lhs (fork46_outs_0),
    .lhs_valid (fork46_outs_0_valid),
    .lhs_ready (fork46_outs_0_ready),
    .rhs (constant508_outs),
    .rhs_valid (constant508_outs_valid),
    .rhs_ready (constant508_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi15_result),
    .result_valid (cmpi15_result_valid),
    .result_ready (cmpi15_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork48(
    .ins (cmpi15_result),
    .ins_valid (cmpi15_result_valid),
    .ins_ready (cmpi15_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork48_outs_8, fork48_outs_7, fork48_outs_6, fork48_outs_5, fork48_outs_4, fork48_outs_3, fork48_outs_2, fork48_outs_1, fork48_outs_0}),
    .outs_valid ({fork48_outs_8_valid, fork48_outs_7_valid, fork48_outs_6_valid, fork48_outs_5_valid, fork48_outs_4_valid, fork48_outs_3_valid, fork48_outs_2_valid, fork48_outs_1_valid, fork48_outs_0_valid}),
    .outs_ready ({fork48_outs_8_ready, fork48_outs_7_ready, fork48_outs_6_ready, fork48_outs_5_ready, fork48_outs_4_ready, fork48_outs_3_ready, fork48_outs_2_ready, fork48_outs_1_ready, fork48_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br167(
    .condition (fork48_outs_5),
    .condition_valid (fork48_outs_5_valid),
    .condition_ready (fork48_outs_5_ready),
    .data (constant328_outs),
    .data_valid (constant328_outs_valid),
    .data_ready (constant328_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br167_trueOut),
    .trueOut_valid (cond_br167_trueOut_valid),
    .trueOut_ready (cond_br167_trueOut_ready),
    .falseOut (cond_br167_falseOut),
    .falseOut_valid (cond_br167_falseOut_valid),
    .falseOut_ready (cond_br167_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink120(
    .ins (cond_br167_falseOut),
    .ins_valid (cond_br167_falseOut_valid),
    .ins_ready (cond_br167_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(31)) cond_br168(
    .condition (fork48_outs_7),
    .condition_valid (fork48_outs_7_valid),
    .condition_ready (fork48_outs_7_ready),
    .data (constant506_outs),
    .data_valid (constant506_outs_valid),
    .data_ready (constant506_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br168_trueOut),
    .trueOut_valid (cond_br168_trueOut_valid),
    .trueOut_ready (cond_br168_trueOut_ready),
    .falseOut (cond_br168_falseOut),
    .falseOut_valid (cond_br168_falseOut_valid),
    .falseOut_ready (cond_br168_falseOut_ready)
  );

  sink #(.DATA_TYPE(31)) sink121(
    .ins (cond_br168_falseOut),
    .ins_valid (cond_br168_falseOut_valid),
    .ins_ready (cond_br168_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(31), .OUTPUT_TYPE(33)) extsi180(
    .ins (cond_br168_trueOut),
    .ins_valid (cond_br168_trueOut_valid),
    .ins_ready (cond_br168_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi180_outs),
    .outs_valid (extsi180_outs_valid),
    .outs_ready (extsi180_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br169(
    .condition (fork48_outs_4),
    .condition_valid (fork48_outs_4_valid),
    .condition_ready (fork48_outs_4_ready),
    .data (constant330_outs),
    .data_valid (constant330_outs_valid),
    .data_ready (constant330_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br169_trueOut),
    .trueOut_valid (cond_br169_trueOut_valid),
    .trueOut_ready (cond_br169_trueOut_ready),
    .falseOut (cond_br169_falseOut),
    .falseOut_valid (cond_br169_falseOut_valid),
    .falseOut_ready (cond_br169_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink122(
    .ins (cond_br169_falseOut),
    .ins_valid (cond_br169_falseOut_valid),
    .ins_ready (cond_br169_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(21)) cond_br170(
    .condition (fork48_outs_6),
    .condition_valid (fork48_outs_6_valid),
    .condition_ready (fork48_outs_6_ready),
    .data (constant507_outs),
    .data_valid (constant507_outs_valid),
    .data_ready (constant507_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br170_trueOut),
    .trueOut_valid (cond_br170_trueOut_valid),
    .trueOut_ready (cond_br170_trueOut_ready),
    .falseOut (cond_br170_falseOut),
    .falseOut_valid (cond_br170_falseOut_valid),
    .falseOut_ready (cond_br170_falseOut_ready)
  );

  sink #(.DATA_TYPE(21)) sink123(
    .ins (cond_br170_falseOut),
    .ins_valid (cond_br170_falseOut_valid),
    .ins_ready (cond_br170_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(21), .OUTPUT_TYPE(22)) extsi181(
    .ins (cond_br170_trueOut),
    .ins_valid (cond_br170_trueOut_valid),
    .ins_ready (cond_br170_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi181_outs),
    .outs_valid (extsi181_outs_valid),
    .outs_ready (extsi181_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br171(
    .condition (fork48_outs_3),
    .condition_valid (fork48_outs_3_valid),
    .condition_ready (fork48_outs_3_ready),
    .data (constant332_outs),
    .data_valid (constant332_outs_valid),
    .data_ready (constant332_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br171_trueOut),
    .trueOut_valid (cond_br171_trueOut_valid),
    .trueOut_ready (cond_br171_trueOut_ready),
    .falseOut (cond_br171_falseOut),
    .falseOut_valid (cond_br171_falseOut_valid),
    .falseOut_ready (cond_br171_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink124(
    .ins (cond_br171_falseOut),
    .ins_valid (cond_br171_falseOut_valid),
    .ins_ready (cond_br171_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br172(
    .condition (fork48_outs_2),
    .condition_valid (fork48_outs_2_valid),
    .condition_ready (fork48_outs_2_ready),
    .data (constant333_outs),
    .data_valid (constant333_outs_valid),
    .data_ready (constant333_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br172_trueOut),
    .trueOut_valid (cond_br172_trueOut_valid),
    .trueOut_ready (cond_br172_trueOut_ready),
    .falseOut (cond_br172_falseOut),
    .falseOut_valid (cond_br172_falseOut_valid),
    .falseOut_ready (cond_br172_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink125(
    .ins (cond_br172_falseOut),
    .ins_valid (cond_br172_falseOut_valid),
    .ins_ready (cond_br172_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer84(
    .ins (cond_br164_falseOut),
    .ins_valid (cond_br164_falseOut_valid),
    .ins_ready (cond_br164_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer84_outs),
    .outs_valid (buffer84_outs_valid),
    .outs_ready (buffer84_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer85(
    .ins (buffer84_outs),
    .ins_valid (buffer84_outs_valid),
    .ins_ready (buffer84_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer85_outs),
    .outs_valid (buffer85_outs_valid),
    .outs_ready (buffer85_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br173(
    .condition (fork48_outs_0),
    .condition_valid (fork48_outs_0_valid),
    .condition_ready (fork48_outs_0_ready),
    .data (buffer85_outs),
    .data_valid (buffer85_outs_valid),
    .data_ready (buffer85_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br173_trueOut),
    .trueOut_valid (cond_br173_trueOut_valid),
    .trueOut_ready (cond_br173_trueOut_ready),
    .falseOut (cond_br173_falseOut),
    .falseOut_valid (cond_br173_falseOut_valid),
    .falseOut_ready (cond_br173_falseOut_ready)
  );

  cond_br_dataless cond_br174(
    .condition (fork48_outs_1),
    .condition_valid (fork48_outs_1_valid),
    .condition_ready (fork48_outs_1_ready),
    .data_valid (fork47_outs_6_valid),
    .data_ready (fork47_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br174_trueOut_valid),
    .trueOut_ready (cond_br174_trueOut_ready),
    .falseOut_valid (cond_br174_falseOut_valid),
    .falseOut_ready (cond_br174_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br175(
    .condition (fork48_outs_8),
    .condition_valid (fork48_outs_8_valid),
    .condition_ready (fork48_outs_8_ready),
    .data (fork46_outs_1),
    .data_valid (fork46_outs_1_valid),
    .data_ready (fork46_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br175_trueOut),
    .trueOut_valid (cond_br175_trueOut_valid),
    .trueOut_ready (cond_br175_trueOut_ready),
    .falseOut (cond_br175_falseOut),
    .falseOut_valid (cond_br175_falseOut_valid),
    .falseOut_ready (cond_br175_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink126(
    .ins (cond_br175_trueOut),
    .ins_valid (cond_br175_trueOut_valid),
    .ins_ready (cond_br175_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer92(
    .ins (cond_br175_falseOut),
    .ins_valid (cond_br175_falseOut_valid),
    .ins_ready (cond_br175_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer92_outs),
    .outs_valid (buffer92_outs_valid),
    .outs_ready (buffer92_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer93(
    .ins (buffer92_outs),
    .ins_valid (buffer92_outs_valid),
    .ins_ready (buffer92_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer93_outs),
    .outs_valid (buffer93_outs_valid),
    .outs_ready (buffer93_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork49(
    .ins (buffer93_outs),
    .ins_valid (buffer93_outs_valid),
    .ins_ready (buffer93_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork49_outs_1, fork49_outs_0}),
    .outs_valid ({fork49_outs_1_valid, fork49_outs_0_valid}),
    .outs_ready ({fork49_outs_1_ready, fork49_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi182(
    .ins (fork49_outs_0),
    .ins_valid (fork49_outs_0_valid),
    .ins_ready (fork49_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi182_outs),
    .outs_valid (extsi182_outs_valid),
    .outs_ready (extsi182_outs_ready)
  );

  oehb_dataless buffer94(
    .ins_valid (cond_br174_falseOut_valid),
    .ins_ready (cond_br174_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer94_outs_valid),
    .outs_ready (buffer94_outs_ready)
  );

  tehb_dataless buffer95(
    .ins_valid (buffer94_outs_valid),
    .ins_ready (buffer94_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer95_outs_valid),
    .outs_ready (buffer95_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork50(
    .ins_valid (buffer95_outs_valid),
    .ins_ready (buffer95_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork50_outs_6_valid, fork50_outs_5_valid, fork50_outs_4_valid, fork50_outs_3_valid, fork50_outs_2_valid, fork50_outs_1_valid, fork50_outs_0_valid}),
    .outs_ready ({fork50_outs_6_ready, fork50_outs_5_ready, fork50_outs_4_ready, fork50_outs_3_ready, fork50_outs_2_ready, fork50_outs_1_ready, fork50_outs_0_ready})
  );

  handshake_constant_112 #(.DATA_WIDTH(37)) constant335(
    .ctrl_valid (fork50_outs_5_valid),
    .ctrl_ready (fork50_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant335_outs),
    .outs_valid (constant335_outs_valid),
    .outs_ready (constant335_outs_ready)
  );

  handshake_constant_113 #(.DATA_WIDTH(30)) constant509(
    .ctrl_valid (fork50_outs_1_valid),
    .ctrl_ready (fork50_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant509_outs),
    .outs_valid (constant509_outs_valid),
    .outs_ready (constant509_outs_ready)
  );

  handshake_constant_114 #(.DATA_WIDTH(27)) constant337(
    .ctrl_valid (fork50_outs_4_valid),
    .ctrl_ready (fork50_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant337_outs),
    .outs_valid (constant337_outs_valid),
    .outs_ready (constant337_outs_ready)
  );

  handshake_constant_115 #(.DATA_WIDTH(20)) constant510(
    .ctrl_valid (fork50_outs_0_valid),
    .ctrl_ready (fork50_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant510_outs),
    .outs_valid (constant510_outs_valid),
    .outs_ready (constant510_outs_ready)
  );

  handshake_constant_116 #(.DATA_WIDTH(17)) constant339(
    .ctrl_valid (fork50_outs_3_valid),
    .ctrl_ready (fork50_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant339_outs),
    .outs_valid (constant339_outs_valid),
    .outs_ready (constant339_outs_ready)
  );

  handshake_constant_117 #(.DATA_WIDTH(12)) constant340(
    .ctrl_valid (fork50_outs_2_valid),
    .ctrl_ready (fork50_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant340_outs),
    .outs_valid (constant340_outs_valid),
    .outs_ready (constant340_outs_ready)
  );

  source source17(
    .clk (clk),
    .rst (rst),
    .outs_valid (source17_outs_valid),
    .outs_ready (source17_outs_ready)
  );

  handshake_constant_118 #(.DATA_WIDTH(6)) constant511(
    .ctrl_valid (source17_outs_valid),
    .ctrl_ready (source17_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant511_outs),
    .outs_valid (constant511_outs_valid),
    .outs_ready (constant511_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi16(
    .lhs (extsi182_outs),
    .lhs_valid (extsi182_outs_valid),
    .lhs_ready (extsi182_outs_ready),
    .rhs (constant511_outs),
    .rhs_valid (constant511_outs_valid),
    .rhs_ready (constant511_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi16_result),
    .result_valid (cmpi16_result_valid),
    .result_ready (cmpi16_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork51(
    .ins (cmpi16_result),
    .ins_valid (cmpi16_result_valid),
    .ins_ready (cmpi16_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork51_outs_8, fork51_outs_7, fork51_outs_6, fork51_outs_5, fork51_outs_4, fork51_outs_3, fork51_outs_2, fork51_outs_1, fork51_outs_0}),
    .outs_valid ({fork51_outs_8_valid, fork51_outs_7_valid, fork51_outs_6_valid, fork51_outs_5_valid, fork51_outs_4_valid, fork51_outs_3_valid, fork51_outs_2_valid, fork51_outs_1_valid, fork51_outs_0_valid}),
    .outs_ready ({fork51_outs_8_ready, fork51_outs_7_ready, fork51_outs_6_ready, fork51_outs_5_ready, fork51_outs_4_ready, fork51_outs_3_ready, fork51_outs_2_ready, fork51_outs_1_ready, fork51_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br176(
    .condition (fork51_outs_5),
    .condition_valid (fork51_outs_5_valid),
    .condition_ready (fork51_outs_5_ready),
    .data (constant335_outs),
    .data_valid (constant335_outs_valid),
    .data_ready (constant335_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br176_trueOut),
    .trueOut_valid (cond_br176_trueOut_valid),
    .trueOut_ready (cond_br176_trueOut_ready),
    .falseOut (cond_br176_falseOut),
    .falseOut_valid (cond_br176_falseOut_valid),
    .falseOut_ready (cond_br176_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink128(
    .ins (cond_br176_falseOut),
    .ins_valid (cond_br176_falseOut_valid),
    .ins_ready (cond_br176_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(30)) cond_br177(
    .condition (fork51_outs_7),
    .condition_valid (fork51_outs_7_valid),
    .condition_ready (fork51_outs_7_ready),
    .data (constant509_outs),
    .data_valid (constant509_outs_valid),
    .data_ready (constant509_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br177_trueOut),
    .trueOut_valid (cond_br177_trueOut_valid),
    .trueOut_ready (cond_br177_trueOut_ready),
    .falseOut (cond_br177_falseOut),
    .falseOut_valid (cond_br177_falseOut_valid),
    .falseOut_ready (cond_br177_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink129(
    .ins (cond_br177_falseOut),
    .ins_valid (cond_br177_falseOut_valid),
    .ins_ready (cond_br177_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(30), .OUTPUT_TYPE(33)) extsi183(
    .ins (cond_br177_trueOut),
    .ins_valid (cond_br177_trueOut_valid),
    .ins_ready (cond_br177_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi183_outs),
    .outs_valid (extsi183_outs_valid),
    .outs_ready (extsi183_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br178(
    .condition (fork51_outs_4),
    .condition_valid (fork51_outs_4_valid),
    .condition_ready (fork51_outs_4_ready),
    .data (constant337_outs),
    .data_valid (constant337_outs_valid),
    .data_ready (constant337_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br178_trueOut),
    .trueOut_valid (cond_br178_trueOut_valid),
    .trueOut_ready (cond_br178_trueOut_ready),
    .falseOut (cond_br178_falseOut),
    .falseOut_valid (cond_br178_falseOut_valid),
    .falseOut_ready (cond_br178_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink130(
    .ins (cond_br178_falseOut),
    .ins_valid (cond_br178_falseOut_valid),
    .ins_ready (cond_br178_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(20)) cond_br179(
    .condition (fork51_outs_6),
    .condition_valid (fork51_outs_6_valid),
    .condition_ready (fork51_outs_6_ready),
    .data (constant510_outs),
    .data_valid (constant510_outs_valid),
    .data_ready (constant510_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br179_trueOut),
    .trueOut_valid (cond_br179_trueOut_valid),
    .trueOut_ready (cond_br179_trueOut_ready),
    .falseOut (cond_br179_falseOut),
    .falseOut_valid (cond_br179_falseOut_valid),
    .falseOut_ready (cond_br179_falseOut_ready)
  );

  sink #(.DATA_TYPE(20)) sink131(
    .ins (cond_br179_falseOut),
    .ins_valid (cond_br179_falseOut_valid),
    .ins_ready (cond_br179_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(20), .OUTPUT_TYPE(22)) extsi184(
    .ins (cond_br179_trueOut),
    .ins_valid (cond_br179_trueOut_valid),
    .ins_ready (cond_br179_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi184_outs),
    .outs_valid (extsi184_outs_valid),
    .outs_ready (extsi184_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br180(
    .condition (fork51_outs_3),
    .condition_valid (fork51_outs_3_valid),
    .condition_ready (fork51_outs_3_ready),
    .data (constant339_outs),
    .data_valid (constant339_outs_valid),
    .data_ready (constant339_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br180_trueOut),
    .trueOut_valid (cond_br180_trueOut_valid),
    .trueOut_ready (cond_br180_trueOut_ready),
    .falseOut (cond_br180_falseOut),
    .falseOut_valid (cond_br180_falseOut_valid),
    .falseOut_ready (cond_br180_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink132(
    .ins (cond_br180_falseOut),
    .ins_valid (cond_br180_falseOut_valid),
    .ins_ready (cond_br180_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(12)) cond_br181(
    .condition (fork51_outs_2),
    .condition_valid (fork51_outs_2_valid),
    .condition_ready (fork51_outs_2_ready),
    .data (constant340_outs),
    .data_valid (constant340_outs_valid),
    .data_ready (constant340_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br181_trueOut),
    .trueOut_valid (cond_br181_trueOut_valid),
    .trueOut_ready (cond_br181_trueOut_ready),
    .falseOut (cond_br181_falseOut),
    .falseOut_valid (cond_br181_falseOut_valid),
    .falseOut_ready (cond_br181_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink133(
    .ins (cond_br181_falseOut),
    .ins_valid (cond_br181_falseOut_valid),
    .ins_ready (cond_br181_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(7)) buffer90(
    .ins (cond_br173_falseOut),
    .ins_valid (cond_br173_falseOut_valid),
    .ins_ready (cond_br173_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer90_outs),
    .outs_valid (buffer90_outs_valid),
    .outs_ready (buffer90_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer91(
    .ins (buffer90_outs),
    .ins_valid (buffer90_outs_valid),
    .ins_ready (buffer90_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer91_outs),
    .outs_valid (buffer91_outs_valid),
    .outs_ready (buffer91_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br182(
    .condition (fork51_outs_0),
    .condition_valid (fork51_outs_0_valid),
    .condition_ready (fork51_outs_0_ready),
    .data (buffer91_outs),
    .data_valid (buffer91_outs_valid),
    .data_ready (buffer91_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br182_trueOut),
    .trueOut_valid (cond_br182_trueOut_valid),
    .trueOut_ready (cond_br182_trueOut_ready),
    .falseOut (cond_br182_falseOut),
    .falseOut_valid (cond_br182_falseOut_valid),
    .falseOut_ready (cond_br182_falseOut_ready)
  );

  cond_br_dataless cond_br183(
    .condition (fork51_outs_1),
    .condition_valid (fork51_outs_1_valid),
    .condition_ready (fork51_outs_1_ready),
    .data_valid (fork50_outs_6_valid),
    .data_ready (fork50_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br183_trueOut_valid),
    .trueOut_ready (cond_br183_trueOut_ready),
    .falseOut_valid (cond_br183_falseOut_valid),
    .falseOut_ready (cond_br183_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br184(
    .condition (fork51_outs_8),
    .condition_valid (fork51_outs_8_valid),
    .condition_ready (fork51_outs_8_ready),
    .data (fork49_outs_1),
    .data_valid (fork49_outs_1_valid),
    .data_ready (fork49_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br184_trueOut),
    .trueOut_valid (cond_br184_trueOut_valid),
    .trueOut_ready (cond_br184_trueOut_ready),
    .falseOut (cond_br184_falseOut),
    .falseOut_valid (cond_br184_falseOut_valid),
    .falseOut_ready (cond_br184_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink134(
    .ins (cond_br184_trueOut),
    .ins_valid (cond_br184_trueOut_valid),
    .ins_ready (cond_br184_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer98(
    .ins (cond_br184_falseOut),
    .ins_valid (cond_br184_falseOut_valid),
    .ins_ready (cond_br184_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer98_outs),
    .outs_valid (buffer98_outs_valid),
    .outs_ready (buffer98_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer99(
    .ins (buffer98_outs),
    .ins_valid (buffer98_outs_valid),
    .ins_ready (buffer98_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer99_outs),
    .outs_valid (buffer99_outs_valid),
    .outs_ready (buffer99_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork52(
    .ins (buffer99_outs),
    .ins_valid (buffer99_outs_valid),
    .ins_ready (buffer99_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork52_outs_1, fork52_outs_0}),
    .outs_valid ({fork52_outs_1_valid, fork52_outs_0_valid}),
    .outs_ready ({fork52_outs_1_ready, fork52_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi185(
    .ins (fork52_outs_0),
    .ins_valid (fork52_outs_0_valid),
    .ins_ready (fork52_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi185_outs),
    .outs_valid (extsi185_outs_valid),
    .outs_ready (extsi185_outs_ready)
  );

  oehb_dataless buffer100(
    .ins_valid (cond_br183_falseOut_valid),
    .ins_ready (cond_br183_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer100_outs_valid),
    .outs_ready (buffer100_outs_ready)
  );

  tehb_dataless buffer101(
    .ins_valid (buffer100_outs_valid),
    .ins_ready (buffer100_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer101_outs_valid),
    .outs_ready (buffer101_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork53(
    .ins_valid (buffer101_outs_valid),
    .ins_ready (buffer101_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork53_outs_6_valid, fork53_outs_5_valid, fork53_outs_4_valid, fork53_outs_3_valid, fork53_outs_2_valid, fork53_outs_1_valid, fork53_outs_0_valid}),
    .outs_ready ({fork53_outs_6_ready, fork53_outs_5_ready, fork53_outs_4_ready, fork53_outs_3_ready, fork53_outs_2_ready, fork53_outs_1_ready, fork53_outs_0_ready})
  );

  handshake_constant_119 #(.DATA_WIDTH(37)) constant342(
    .ctrl_valid (fork53_outs_5_valid),
    .ctrl_ready (fork53_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant342_outs),
    .outs_valid (constant342_outs_valid),
    .outs_ready (constant342_outs_ready)
  );

  handshake_constant_120 #(.DATA_WIDTH(30)) constant512(
    .ctrl_valid (fork53_outs_2_valid),
    .ctrl_ready (fork53_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant512_outs),
    .outs_valid (constant512_outs_valid),
    .outs_ready (constant512_outs_ready)
  );

  handshake_constant_121 #(.DATA_WIDTH(27)) constant344(
    .ctrl_valid (fork53_outs_4_valid),
    .ctrl_ready (fork53_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant344_outs),
    .outs_valid (constant344_outs_valid),
    .outs_ready (constant344_outs_ready)
  );

  handshake_constant_122 #(.DATA_WIDTH(20)) constant513(
    .ctrl_valid (fork53_outs_1_valid),
    .ctrl_ready (fork53_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant513_outs),
    .outs_valid (constant513_outs_valid),
    .outs_ready (constant513_outs_ready)
  );

  handshake_constant_123 #(.DATA_WIDTH(17)) constant346(
    .ctrl_valid (fork53_outs_3_valid),
    .ctrl_ready (fork53_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant346_outs),
    .outs_valid (constant346_outs_valid),
    .outs_ready (constant346_outs_ready)
  );

  handshake_constant_124 #(.DATA_WIDTH(6)) constant514(
    .ctrl_valid (fork53_outs_0_valid),
    .ctrl_ready (fork53_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant514_outs),
    .outs_valid (constant514_outs_valid),
    .outs_ready (constant514_outs_ready)
  );

  source source18(
    .clk (clk),
    .rst (rst),
    .outs_valid (source18_outs_valid),
    .outs_ready (source18_outs_ready)
  );

  handshake_constant_125 #(.DATA_WIDTH(6)) constant515(
    .ctrl_valid (source18_outs_valid),
    .ctrl_ready (source18_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant515_outs),
    .outs_valid (constant515_outs_valid),
    .outs_ready (constant515_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi17(
    .lhs (extsi185_outs),
    .lhs_valid (extsi185_outs_valid),
    .lhs_ready (extsi185_outs_ready),
    .rhs (constant515_outs),
    .rhs_valid (constant515_outs_valid),
    .rhs_ready (constant515_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi17_result),
    .result_valid (cmpi17_result_valid),
    .result_ready (cmpi17_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork54(
    .ins (cmpi17_result),
    .ins_valid (cmpi17_result_valid),
    .ins_ready (cmpi17_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork54_outs_8, fork54_outs_7, fork54_outs_6, fork54_outs_5, fork54_outs_4, fork54_outs_3, fork54_outs_2, fork54_outs_1, fork54_outs_0}),
    .outs_valid ({fork54_outs_8_valid, fork54_outs_7_valid, fork54_outs_6_valid, fork54_outs_5_valid, fork54_outs_4_valid, fork54_outs_3_valid, fork54_outs_2_valid, fork54_outs_1_valid, fork54_outs_0_valid}),
    .outs_ready ({fork54_outs_8_ready, fork54_outs_7_ready, fork54_outs_6_ready, fork54_outs_5_ready, fork54_outs_4_ready, fork54_outs_3_ready, fork54_outs_2_ready, fork54_outs_1_ready, fork54_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br185(
    .condition (fork54_outs_4),
    .condition_valid (fork54_outs_4_valid),
    .condition_ready (fork54_outs_4_ready),
    .data (constant342_outs),
    .data_valid (constant342_outs_valid),
    .data_ready (constant342_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br185_trueOut),
    .trueOut_valid (cond_br185_trueOut_valid),
    .trueOut_ready (cond_br185_trueOut_ready),
    .falseOut (cond_br185_falseOut),
    .falseOut_valid (cond_br185_falseOut_valid),
    .falseOut_ready (cond_br185_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink136(
    .ins (cond_br185_falseOut),
    .ins_valid (cond_br185_falseOut_valid),
    .ins_ready (cond_br185_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(30)) cond_br186(
    .condition (fork54_outs_7),
    .condition_valid (fork54_outs_7_valid),
    .condition_ready (fork54_outs_7_ready),
    .data (constant512_outs),
    .data_valid (constant512_outs_valid),
    .data_ready (constant512_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br186_trueOut),
    .trueOut_valid (cond_br186_trueOut_valid),
    .trueOut_ready (cond_br186_trueOut_ready),
    .falseOut (cond_br186_falseOut),
    .falseOut_valid (cond_br186_falseOut_valid),
    .falseOut_ready (cond_br186_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink137(
    .ins (cond_br186_falseOut),
    .ins_valid (cond_br186_falseOut_valid),
    .ins_ready (cond_br186_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(30), .OUTPUT_TYPE(33)) extsi186(
    .ins (cond_br186_trueOut),
    .ins_valid (cond_br186_trueOut_valid),
    .ins_ready (cond_br186_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi186_outs),
    .outs_valid (extsi186_outs_valid),
    .outs_ready (extsi186_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br187(
    .condition (fork54_outs_3),
    .condition_valid (fork54_outs_3_valid),
    .condition_ready (fork54_outs_3_ready),
    .data (constant344_outs),
    .data_valid (constant344_outs_valid),
    .data_ready (constant344_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br187_trueOut),
    .trueOut_valid (cond_br187_trueOut_valid),
    .trueOut_ready (cond_br187_trueOut_ready),
    .falseOut (cond_br187_falseOut),
    .falseOut_valid (cond_br187_falseOut_valid),
    .falseOut_ready (cond_br187_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink138(
    .ins (cond_br187_falseOut),
    .ins_valid (cond_br187_falseOut_valid),
    .ins_ready (cond_br187_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(20)) cond_br188(
    .condition (fork54_outs_6),
    .condition_valid (fork54_outs_6_valid),
    .condition_ready (fork54_outs_6_ready),
    .data (constant513_outs),
    .data_valid (constant513_outs_valid),
    .data_ready (constant513_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br188_trueOut),
    .trueOut_valid (cond_br188_trueOut_valid),
    .trueOut_ready (cond_br188_trueOut_ready),
    .falseOut (cond_br188_falseOut),
    .falseOut_valid (cond_br188_falseOut_valid),
    .falseOut_ready (cond_br188_falseOut_ready)
  );

  sink #(.DATA_TYPE(20)) sink139(
    .ins (cond_br188_falseOut),
    .ins_valid (cond_br188_falseOut_valid),
    .ins_ready (cond_br188_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(20), .OUTPUT_TYPE(22)) extsi187(
    .ins (cond_br188_trueOut),
    .ins_valid (cond_br188_trueOut_valid),
    .ins_ready (cond_br188_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi187_outs),
    .outs_valid (extsi187_outs_valid),
    .outs_ready (extsi187_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br189(
    .condition (fork54_outs_2),
    .condition_valid (fork54_outs_2_valid),
    .condition_ready (fork54_outs_2_ready),
    .data (constant346_outs),
    .data_valid (constant346_outs_valid),
    .data_ready (constant346_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br189_trueOut),
    .trueOut_valid (cond_br189_trueOut_valid),
    .trueOut_ready (cond_br189_trueOut_ready),
    .falseOut (cond_br189_falseOut),
    .falseOut_valid (cond_br189_falseOut_valid),
    .falseOut_ready (cond_br189_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink140(
    .ins (cond_br189_falseOut),
    .ins_valid (cond_br189_falseOut_valid),
    .ins_ready (cond_br189_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(6)) cond_br190(
    .condition (fork54_outs_5),
    .condition_valid (fork54_outs_5_valid),
    .condition_ready (fork54_outs_5_ready),
    .data (constant514_outs),
    .data_valid (constant514_outs_valid),
    .data_ready (constant514_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br190_trueOut),
    .trueOut_valid (cond_br190_trueOut_valid),
    .trueOut_ready (cond_br190_trueOut_ready),
    .falseOut (cond_br190_falseOut),
    .falseOut_valid (cond_br190_falseOut_valid),
    .falseOut_ready (cond_br190_falseOut_ready)
  );

  sink #(.DATA_TYPE(6)) sink141(
    .ins (cond_br190_falseOut),
    .ins_valid (cond_br190_falseOut_valid),
    .ins_ready (cond_br190_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(12)) extsi188(
    .ins (cond_br190_trueOut),
    .ins_valid (cond_br190_trueOut_valid),
    .ins_ready (cond_br190_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi188_outs),
    .outs_valid (extsi188_outs_valid),
    .outs_ready (extsi188_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer96(
    .ins (cond_br182_falseOut),
    .ins_valid (cond_br182_falseOut_valid),
    .ins_ready (cond_br182_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer96_outs),
    .outs_valid (buffer96_outs_valid),
    .outs_ready (buffer96_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer97(
    .ins (buffer96_outs),
    .ins_valid (buffer96_outs_valid),
    .ins_ready (buffer96_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer97_outs),
    .outs_valid (buffer97_outs_valid),
    .outs_ready (buffer97_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br191(
    .condition (fork54_outs_0),
    .condition_valid (fork54_outs_0_valid),
    .condition_ready (fork54_outs_0_ready),
    .data (buffer97_outs),
    .data_valid (buffer97_outs_valid),
    .data_ready (buffer97_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br191_trueOut),
    .trueOut_valid (cond_br191_trueOut_valid),
    .trueOut_ready (cond_br191_trueOut_ready),
    .falseOut (cond_br191_falseOut),
    .falseOut_valid (cond_br191_falseOut_valid),
    .falseOut_ready (cond_br191_falseOut_ready)
  );

  cond_br_dataless cond_br192(
    .condition (fork54_outs_1),
    .condition_valid (fork54_outs_1_valid),
    .condition_ready (fork54_outs_1_ready),
    .data_valid (fork53_outs_6_valid),
    .data_ready (fork53_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br192_trueOut_valid),
    .trueOut_ready (cond_br192_trueOut_ready),
    .falseOut_valid (cond_br192_falseOut_valid),
    .falseOut_ready (cond_br192_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br193(
    .condition (fork54_outs_8),
    .condition_valid (fork54_outs_8_valid),
    .condition_ready (fork54_outs_8_ready),
    .data (fork52_outs_1),
    .data_valid (fork52_outs_1_valid),
    .data_ready (fork52_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br193_trueOut),
    .trueOut_valid (cond_br193_trueOut_valid),
    .trueOut_ready (cond_br193_trueOut_ready),
    .falseOut (cond_br193_falseOut),
    .falseOut_valid (cond_br193_falseOut_valid),
    .falseOut_ready (cond_br193_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink142(
    .ins (cond_br193_trueOut),
    .ins_valid (cond_br193_trueOut_valid),
    .ins_ready (cond_br193_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer104(
    .ins (cond_br193_falseOut),
    .ins_valid (cond_br193_falseOut_valid),
    .ins_ready (cond_br193_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer104_outs),
    .outs_valid (buffer104_outs_valid),
    .outs_ready (buffer104_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer105(
    .ins (buffer104_outs),
    .ins_valid (buffer104_outs_valid),
    .ins_ready (buffer104_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer105_outs),
    .outs_valid (buffer105_outs_valid),
    .outs_ready (buffer105_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork55(
    .ins (buffer105_outs),
    .ins_valid (buffer105_outs_valid),
    .ins_ready (buffer105_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork55_outs_1, fork55_outs_0}),
    .outs_valid ({fork55_outs_1_valid, fork55_outs_0_valid}),
    .outs_ready ({fork55_outs_1_ready, fork55_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi189(
    .ins (fork55_outs_0),
    .ins_valid (fork55_outs_0_valid),
    .ins_ready (fork55_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi189_outs),
    .outs_valid (extsi189_outs_valid),
    .outs_ready (extsi189_outs_ready)
  );

  oehb_dataless buffer106(
    .ins_valid (cond_br192_falseOut_valid),
    .ins_ready (cond_br192_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer106_outs_valid),
    .outs_ready (buffer106_outs_ready)
  );

  tehb_dataless buffer107(
    .ins_valid (buffer106_outs_valid),
    .ins_ready (buffer106_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer107_outs_valid),
    .outs_ready (buffer107_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork56(
    .ins_valid (buffer107_outs_valid),
    .ins_ready (buffer107_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork56_outs_6_valid, fork56_outs_5_valid, fork56_outs_4_valid, fork56_outs_3_valid, fork56_outs_2_valid, fork56_outs_1_valid, fork56_outs_0_valid}),
    .outs_ready ({fork56_outs_6_ready, fork56_outs_5_ready, fork56_outs_4_ready, fork56_outs_3_ready, fork56_outs_2_ready, fork56_outs_1_ready, fork56_outs_0_ready})
  );

  handshake_constant_126 #(.DATA_WIDTH(37)) constant349(
    .ctrl_valid (fork56_outs_5_valid),
    .ctrl_ready (fork56_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant349_outs),
    .outs_valid (constant349_outs_valid),
    .outs_ready (constant349_outs_ready)
  );

  handshake_constant_127 #(.DATA_WIDTH(30)) constant516(
    .ctrl_valid (fork56_outs_2_valid),
    .ctrl_ready (fork56_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant516_outs),
    .outs_valid (constant516_outs_valid),
    .outs_ready (constant516_outs_ready)
  );

  handshake_constant_128 #(.DATA_WIDTH(27)) constant351(
    .ctrl_valid (fork56_outs_4_valid),
    .ctrl_ready (fork56_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant351_outs),
    .outs_valid (constant351_outs_valid),
    .outs_ready (constant351_outs_ready)
  );

  handshake_constant_129 #(.DATA_WIDTH(20)) constant517(
    .ctrl_valid (fork56_outs_1_valid),
    .ctrl_ready (fork56_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant517_outs),
    .outs_valid (constant517_outs_valid),
    .outs_ready (constant517_outs_ready)
  );

  handshake_constant_130 #(.DATA_WIDTH(17)) constant353(
    .ctrl_valid (fork56_outs_3_valid),
    .ctrl_ready (fork56_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant353_outs),
    .outs_valid (constant353_outs_valid),
    .outs_ready (constant353_outs_ready)
  );

  handshake_constant_131 #(.DATA_WIDTH(7)) constant518(
    .ctrl_valid (fork56_outs_0_valid),
    .ctrl_ready (fork56_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant518_outs),
    .outs_valid (constant518_outs_valid),
    .outs_ready (constant518_outs_ready)
  );

  source source19(
    .clk (clk),
    .rst (rst),
    .outs_valid (source19_outs_valid),
    .outs_ready (source19_outs_ready)
  );

  handshake_constant_132 #(.DATA_WIDTH(6)) constant519(
    .ctrl_valid (source19_outs_valid),
    .ctrl_ready (source19_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant519_outs),
    .outs_valid (constant519_outs_valid),
    .outs_ready (constant519_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi18(
    .lhs (extsi189_outs),
    .lhs_valid (extsi189_outs_valid),
    .lhs_ready (extsi189_outs_ready),
    .rhs (constant519_outs),
    .rhs_valid (constant519_outs_valid),
    .rhs_ready (constant519_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi18_result),
    .result_valid (cmpi18_result_valid),
    .result_ready (cmpi18_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork57(
    .ins (cmpi18_result),
    .ins_valid (cmpi18_result_valid),
    .ins_ready (cmpi18_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork57_outs_8, fork57_outs_7, fork57_outs_6, fork57_outs_5, fork57_outs_4, fork57_outs_3, fork57_outs_2, fork57_outs_1, fork57_outs_0}),
    .outs_valid ({fork57_outs_8_valid, fork57_outs_7_valid, fork57_outs_6_valid, fork57_outs_5_valid, fork57_outs_4_valid, fork57_outs_3_valid, fork57_outs_2_valid, fork57_outs_1_valid, fork57_outs_0_valid}),
    .outs_ready ({fork57_outs_8_ready, fork57_outs_7_ready, fork57_outs_6_ready, fork57_outs_5_ready, fork57_outs_4_ready, fork57_outs_3_ready, fork57_outs_2_ready, fork57_outs_1_ready, fork57_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br194(
    .condition (fork57_outs_4),
    .condition_valid (fork57_outs_4_valid),
    .condition_ready (fork57_outs_4_ready),
    .data (constant349_outs),
    .data_valid (constant349_outs_valid),
    .data_ready (constant349_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br194_trueOut),
    .trueOut_valid (cond_br194_trueOut_valid),
    .trueOut_ready (cond_br194_trueOut_ready),
    .falseOut (cond_br194_falseOut),
    .falseOut_valid (cond_br194_falseOut_valid),
    .falseOut_ready (cond_br194_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink144(
    .ins (cond_br194_falseOut),
    .ins_valid (cond_br194_falseOut_valid),
    .ins_ready (cond_br194_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(30)) cond_br195(
    .condition (fork57_outs_7),
    .condition_valid (fork57_outs_7_valid),
    .condition_ready (fork57_outs_7_ready),
    .data (constant516_outs),
    .data_valid (constant516_outs_valid),
    .data_ready (constant516_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br195_trueOut),
    .trueOut_valid (cond_br195_trueOut_valid),
    .trueOut_ready (cond_br195_trueOut_ready),
    .falseOut (cond_br195_falseOut),
    .falseOut_valid (cond_br195_falseOut_valid),
    .falseOut_ready (cond_br195_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink145(
    .ins (cond_br195_falseOut),
    .ins_valid (cond_br195_falseOut_valid),
    .ins_ready (cond_br195_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(30), .OUTPUT_TYPE(33)) extsi190(
    .ins (cond_br195_trueOut),
    .ins_valid (cond_br195_trueOut_valid),
    .ins_ready (cond_br195_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi190_outs),
    .outs_valid (extsi190_outs_valid),
    .outs_ready (extsi190_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br196(
    .condition (fork57_outs_3),
    .condition_valid (fork57_outs_3_valid),
    .condition_ready (fork57_outs_3_ready),
    .data (constant351_outs),
    .data_valid (constant351_outs_valid),
    .data_ready (constant351_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br196_trueOut),
    .trueOut_valid (cond_br196_trueOut_valid),
    .trueOut_ready (cond_br196_trueOut_ready),
    .falseOut (cond_br196_falseOut),
    .falseOut_valid (cond_br196_falseOut_valid),
    .falseOut_ready (cond_br196_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink146(
    .ins (cond_br196_falseOut),
    .ins_valid (cond_br196_falseOut_valid),
    .ins_ready (cond_br196_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(20)) cond_br197(
    .condition (fork57_outs_6),
    .condition_valid (fork57_outs_6_valid),
    .condition_ready (fork57_outs_6_ready),
    .data (constant517_outs),
    .data_valid (constant517_outs_valid),
    .data_ready (constant517_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br197_trueOut),
    .trueOut_valid (cond_br197_trueOut_valid),
    .trueOut_ready (cond_br197_trueOut_ready),
    .falseOut (cond_br197_falseOut),
    .falseOut_valid (cond_br197_falseOut_valid),
    .falseOut_ready (cond_br197_falseOut_ready)
  );

  sink #(.DATA_TYPE(20)) sink147(
    .ins (cond_br197_falseOut),
    .ins_valid (cond_br197_falseOut_valid),
    .ins_ready (cond_br197_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(20), .OUTPUT_TYPE(22)) extsi191(
    .ins (cond_br197_trueOut),
    .ins_valid (cond_br197_trueOut_valid),
    .ins_ready (cond_br197_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi191_outs),
    .outs_valid (extsi191_outs_valid),
    .outs_ready (extsi191_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br198(
    .condition (fork57_outs_2),
    .condition_valid (fork57_outs_2_valid),
    .condition_ready (fork57_outs_2_ready),
    .data (constant353_outs),
    .data_valid (constant353_outs_valid),
    .data_ready (constant353_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br198_trueOut),
    .trueOut_valid (cond_br198_trueOut_valid),
    .trueOut_ready (cond_br198_trueOut_ready),
    .falseOut (cond_br198_falseOut),
    .falseOut_valid (cond_br198_falseOut_valid),
    .falseOut_ready (cond_br198_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink148(
    .ins (cond_br198_falseOut),
    .ins_valid (cond_br198_falseOut_valid),
    .ins_ready (cond_br198_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br199(
    .condition (fork57_outs_5),
    .condition_valid (fork57_outs_5_valid),
    .condition_ready (fork57_outs_5_ready),
    .data (constant518_outs),
    .data_valid (constant518_outs_valid),
    .data_ready (constant518_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br199_trueOut),
    .trueOut_valid (cond_br199_trueOut_valid),
    .trueOut_ready (cond_br199_trueOut_ready),
    .falseOut (cond_br199_falseOut),
    .falseOut_valid (cond_br199_falseOut_valid),
    .falseOut_ready (cond_br199_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink149(
    .ins (cond_br199_falseOut),
    .ins_valid (cond_br199_falseOut_valid),
    .ins_ready (cond_br199_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(12)) extsi192(
    .ins (cond_br199_trueOut),
    .ins_valid (cond_br199_trueOut_valid),
    .ins_ready (cond_br199_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi192_outs),
    .outs_valid (extsi192_outs_valid),
    .outs_ready (extsi192_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer102(
    .ins (cond_br191_falseOut),
    .ins_valid (cond_br191_falseOut_valid),
    .ins_ready (cond_br191_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer102_outs),
    .outs_valid (buffer102_outs_valid),
    .outs_ready (buffer102_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer103(
    .ins (buffer102_outs),
    .ins_valid (buffer102_outs_valid),
    .ins_ready (buffer102_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer103_outs),
    .outs_valid (buffer103_outs_valid),
    .outs_ready (buffer103_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br200(
    .condition (fork57_outs_0),
    .condition_valid (fork57_outs_0_valid),
    .condition_ready (fork57_outs_0_ready),
    .data (buffer103_outs),
    .data_valid (buffer103_outs_valid),
    .data_ready (buffer103_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br200_trueOut),
    .trueOut_valid (cond_br200_trueOut_valid),
    .trueOut_ready (cond_br200_trueOut_ready),
    .falseOut (cond_br200_falseOut),
    .falseOut_valid (cond_br200_falseOut_valid),
    .falseOut_ready (cond_br200_falseOut_ready)
  );

  cond_br_dataless cond_br201(
    .condition (fork57_outs_1),
    .condition_valid (fork57_outs_1_valid),
    .condition_ready (fork57_outs_1_ready),
    .data_valid (fork56_outs_6_valid),
    .data_ready (fork56_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br201_trueOut_valid),
    .trueOut_ready (cond_br201_trueOut_ready),
    .falseOut_valid (cond_br201_falseOut_valid),
    .falseOut_ready (cond_br201_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br202(
    .condition (fork57_outs_8),
    .condition_valid (fork57_outs_8_valid),
    .condition_ready (fork57_outs_8_ready),
    .data (fork55_outs_1),
    .data_valid (fork55_outs_1_valid),
    .data_ready (fork55_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br202_trueOut),
    .trueOut_valid (cond_br202_trueOut_valid),
    .trueOut_ready (cond_br202_trueOut_ready),
    .falseOut (cond_br202_falseOut),
    .falseOut_valid (cond_br202_falseOut_valid),
    .falseOut_ready (cond_br202_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink150(
    .ins (cond_br202_trueOut),
    .ins_valid (cond_br202_trueOut_valid),
    .ins_ready (cond_br202_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer110(
    .ins (cond_br202_falseOut),
    .ins_valid (cond_br202_falseOut_valid),
    .ins_ready (cond_br202_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer110_outs),
    .outs_valid (buffer110_outs_valid),
    .outs_ready (buffer110_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer111(
    .ins (buffer110_outs),
    .ins_valid (buffer110_outs_valid),
    .ins_ready (buffer110_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer111_outs),
    .outs_valid (buffer111_outs_valid),
    .outs_ready (buffer111_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork58(
    .ins (buffer111_outs),
    .ins_valid (buffer111_outs_valid),
    .ins_ready (buffer111_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork58_outs_1, fork58_outs_0}),
    .outs_valid ({fork58_outs_1_valid, fork58_outs_0_valid}),
    .outs_ready ({fork58_outs_1_ready, fork58_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi193(
    .ins (fork58_outs_0),
    .ins_valid (fork58_outs_0_valid),
    .ins_ready (fork58_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi193_outs),
    .outs_valid (extsi193_outs_valid),
    .outs_ready (extsi193_outs_ready)
  );

  oehb_dataless buffer112(
    .ins_valid (cond_br201_falseOut_valid),
    .ins_ready (cond_br201_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer112_outs_valid),
    .outs_ready (buffer112_outs_ready)
  );

  tehb_dataless buffer113(
    .ins_valid (buffer112_outs_valid),
    .ins_ready (buffer112_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer113_outs_valid),
    .outs_ready (buffer113_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork59(
    .ins_valid (buffer113_outs_valid),
    .ins_ready (buffer113_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork59_outs_6_valid, fork59_outs_5_valid, fork59_outs_4_valid, fork59_outs_3_valid, fork59_outs_2_valid, fork59_outs_1_valid, fork59_outs_0_valid}),
    .outs_ready ({fork59_outs_6_ready, fork59_outs_5_ready, fork59_outs_4_ready, fork59_outs_3_ready, fork59_outs_2_ready, fork59_outs_1_ready, fork59_outs_0_ready})
  );

  handshake_constant_133 #(.DATA_WIDTH(37)) constant356(
    .ctrl_valid (fork59_outs_5_valid),
    .ctrl_ready (fork59_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant356_outs),
    .outs_valid (constant356_outs_valid),
    .outs_ready (constant356_outs_ready)
  );

  handshake_constant_134 #(.DATA_WIDTH(30)) constant520(
    .ctrl_valid (fork59_outs_2_valid),
    .ctrl_ready (fork59_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant520_outs),
    .outs_valid (constant520_outs_valid),
    .outs_ready (constant520_outs_ready)
  );

  handshake_constant_135 #(.DATA_WIDTH(27)) constant358(
    .ctrl_valid (fork59_outs_4_valid),
    .ctrl_ready (fork59_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant358_outs),
    .outs_valid (constant358_outs_valid),
    .outs_ready (constant358_outs_ready)
  );

  handshake_constant_136 #(.DATA_WIDTH(20)) constant521(
    .ctrl_valid (fork59_outs_1_valid),
    .ctrl_ready (fork59_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant521_outs),
    .outs_valid (constant521_outs_valid),
    .outs_ready (constant521_outs_ready)
  );

  handshake_constant_137 #(.DATA_WIDTH(17)) constant360(
    .ctrl_valid (fork59_outs_3_valid),
    .ctrl_ready (fork59_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant360_outs),
    .outs_valid (constant360_outs_valid),
    .outs_ready (constant360_outs_ready)
  );

  handshake_constant_138 #(.DATA_WIDTH(7)) constant522(
    .ctrl_valid (fork59_outs_0_valid),
    .ctrl_ready (fork59_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant522_outs),
    .outs_valid (constant522_outs_valid),
    .outs_ready (constant522_outs_ready)
  );

  source source20(
    .clk (clk),
    .rst (rst),
    .outs_valid (source20_outs_valid),
    .outs_ready (source20_outs_ready)
  );

  handshake_constant_139 #(.DATA_WIDTH(6)) constant523(
    .ctrl_valid (source20_outs_valid),
    .ctrl_ready (source20_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant523_outs),
    .outs_valid (constant523_outs_valid),
    .outs_ready (constant523_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi19(
    .lhs (extsi193_outs),
    .lhs_valid (extsi193_outs_valid),
    .lhs_ready (extsi193_outs_ready),
    .rhs (constant523_outs),
    .rhs_valid (constant523_outs_valid),
    .rhs_ready (constant523_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi19_result),
    .result_valid (cmpi19_result_valid),
    .result_ready (cmpi19_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork60(
    .ins (cmpi19_result),
    .ins_valid (cmpi19_result_valid),
    .ins_ready (cmpi19_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork60_outs_8, fork60_outs_7, fork60_outs_6, fork60_outs_5, fork60_outs_4, fork60_outs_3, fork60_outs_2, fork60_outs_1, fork60_outs_0}),
    .outs_valid ({fork60_outs_8_valid, fork60_outs_7_valid, fork60_outs_6_valid, fork60_outs_5_valid, fork60_outs_4_valid, fork60_outs_3_valid, fork60_outs_2_valid, fork60_outs_1_valid, fork60_outs_0_valid}),
    .outs_ready ({fork60_outs_8_ready, fork60_outs_7_ready, fork60_outs_6_ready, fork60_outs_5_ready, fork60_outs_4_ready, fork60_outs_3_ready, fork60_outs_2_ready, fork60_outs_1_ready, fork60_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br203(
    .condition (fork60_outs_4),
    .condition_valid (fork60_outs_4_valid),
    .condition_ready (fork60_outs_4_ready),
    .data (constant356_outs),
    .data_valid (constant356_outs_valid),
    .data_ready (constant356_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br203_trueOut),
    .trueOut_valid (cond_br203_trueOut_valid),
    .trueOut_ready (cond_br203_trueOut_ready),
    .falseOut (cond_br203_falseOut),
    .falseOut_valid (cond_br203_falseOut_valid),
    .falseOut_ready (cond_br203_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink152(
    .ins (cond_br203_falseOut),
    .ins_valid (cond_br203_falseOut_valid),
    .ins_ready (cond_br203_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(30)) cond_br204(
    .condition (fork60_outs_7),
    .condition_valid (fork60_outs_7_valid),
    .condition_ready (fork60_outs_7_ready),
    .data (constant520_outs),
    .data_valid (constant520_outs_valid),
    .data_ready (constant520_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br204_trueOut),
    .trueOut_valid (cond_br204_trueOut_valid),
    .trueOut_ready (cond_br204_trueOut_ready),
    .falseOut (cond_br204_falseOut),
    .falseOut_valid (cond_br204_falseOut_valid),
    .falseOut_ready (cond_br204_falseOut_ready)
  );

  sink #(.DATA_TYPE(30)) sink153(
    .ins (cond_br204_falseOut),
    .ins_valid (cond_br204_falseOut_valid),
    .ins_ready (cond_br204_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(30), .OUTPUT_TYPE(33)) extsi194(
    .ins (cond_br204_trueOut),
    .ins_valid (cond_br204_trueOut_valid),
    .ins_ready (cond_br204_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi194_outs),
    .outs_valid (extsi194_outs_valid),
    .outs_ready (extsi194_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br205(
    .condition (fork60_outs_3),
    .condition_valid (fork60_outs_3_valid),
    .condition_ready (fork60_outs_3_ready),
    .data (constant358_outs),
    .data_valid (constant358_outs_valid),
    .data_ready (constant358_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br205_trueOut),
    .trueOut_valid (cond_br205_trueOut_valid),
    .trueOut_ready (cond_br205_trueOut_ready),
    .falseOut (cond_br205_falseOut),
    .falseOut_valid (cond_br205_falseOut_valid),
    .falseOut_ready (cond_br205_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink154(
    .ins (cond_br205_falseOut),
    .ins_valid (cond_br205_falseOut_valid),
    .ins_ready (cond_br205_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(20)) cond_br206(
    .condition (fork60_outs_6),
    .condition_valid (fork60_outs_6_valid),
    .condition_ready (fork60_outs_6_ready),
    .data (constant521_outs),
    .data_valid (constant521_outs_valid),
    .data_ready (constant521_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br206_trueOut),
    .trueOut_valid (cond_br206_trueOut_valid),
    .trueOut_ready (cond_br206_trueOut_ready),
    .falseOut (cond_br206_falseOut),
    .falseOut_valid (cond_br206_falseOut_valid),
    .falseOut_ready (cond_br206_falseOut_ready)
  );

  sink #(.DATA_TYPE(20)) sink155(
    .ins (cond_br206_falseOut),
    .ins_valid (cond_br206_falseOut_valid),
    .ins_ready (cond_br206_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(20), .OUTPUT_TYPE(22)) extsi195(
    .ins (cond_br206_trueOut),
    .ins_valid (cond_br206_trueOut_valid),
    .ins_ready (cond_br206_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi195_outs),
    .outs_valid (extsi195_outs_valid),
    .outs_ready (extsi195_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br207(
    .condition (fork60_outs_2),
    .condition_valid (fork60_outs_2_valid),
    .condition_ready (fork60_outs_2_ready),
    .data (constant360_outs),
    .data_valid (constant360_outs_valid),
    .data_ready (constant360_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br207_trueOut),
    .trueOut_valid (cond_br207_trueOut_valid),
    .trueOut_ready (cond_br207_trueOut_ready),
    .falseOut (cond_br207_falseOut),
    .falseOut_valid (cond_br207_falseOut_valid),
    .falseOut_ready (cond_br207_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink156(
    .ins (cond_br207_falseOut),
    .ins_valid (cond_br207_falseOut_valid),
    .ins_ready (cond_br207_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br208(
    .condition (fork60_outs_5),
    .condition_valid (fork60_outs_5_valid),
    .condition_ready (fork60_outs_5_ready),
    .data (constant522_outs),
    .data_valid (constant522_outs_valid),
    .data_ready (constant522_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br208_trueOut),
    .trueOut_valid (cond_br208_trueOut_valid),
    .trueOut_ready (cond_br208_trueOut_ready),
    .falseOut (cond_br208_falseOut),
    .falseOut_valid (cond_br208_falseOut_valid),
    .falseOut_ready (cond_br208_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink157(
    .ins (cond_br208_falseOut),
    .ins_valid (cond_br208_falseOut_valid),
    .ins_ready (cond_br208_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(12)) extsi196(
    .ins (cond_br208_trueOut),
    .ins_valid (cond_br208_trueOut_valid),
    .ins_ready (cond_br208_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi196_outs),
    .outs_valid (extsi196_outs_valid),
    .outs_ready (extsi196_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer108(
    .ins (cond_br200_falseOut),
    .ins_valid (cond_br200_falseOut_valid),
    .ins_ready (cond_br200_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer108_outs),
    .outs_valid (buffer108_outs_valid),
    .outs_ready (buffer108_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer109(
    .ins (buffer108_outs),
    .ins_valid (buffer108_outs_valid),
    .ins_ready (buffer108_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer109_outs),
    .outs_valid (buffer109_outs_valid),
    .outs_ready (buffer109_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br209(
    .condition (fork60_outs_0),
    .condition_valid (fork60_outs_0_valid),
    .condition_ready (fork60_outs_0_ready),
    .data (buffer109_outs),
    .data_valid (buffer109_outs_valid),
    .data_ready (buffer109_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br209_trueOut),
    .trueOut_valid (cond_br209_trueOut_valid),
    .trueOut_ready (cond_br209_trueOut_ready),
    .falseOut (cond_br209_falseOut),
    .falseOut_valid (cond_br209_falseOut_valid),
    .falseOut_ready (cond_br209_falseOut_ready)
  );

  cond_br_dataless cond_br210(
    .condition (fork60_outs_1),
    .condition_valid (fork60_outs_1_valid),
    .condition_ready (fork60_outs_1_ready),
    .data_valid (fork59_outs_6_valid),
    .data_ready (fork59_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br210_trueOut_valid),
    .trueOut_ready (cond_br210_trueOut_ready),
    .falseOut_valid (cond_br210_falseOut_valid),
    .falseOut_ready (cond_br210_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br211(
    .condition (fork60_outs_8),
    .condition_valid (fork60_outs_8_valid),
    .condition_ready (fork60_outs_8_ready),
    .data (fork58_outs_1),
    .data_valid (fork58_outs_1_valid),
    .data_ready (fork58_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br211_trueOut),
    .trueOut_valid (cond_br211_trueOut_valid),
    .trueOut_ready (cond_br211_trueOut_ready),
    .falseOut (cond_br211_falseOut),
    .falseOut_valid (cond_br211_falseOut_valid),
    .falseOut_ready (cond_br211_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink158(
    .ins (cond_br211_trueOut),
    .ins_valid (cond_br211_trueOut_valid),
    .ins_ready (cond_br211_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer116(
    .ins (cond_br211_falseOut),
    .ins_valid (cond_br211_falseOut_valid),
    .ins_ready (cond_br211_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer116_outs),
    .outs_valid (buffer116_outs_valid),
    .outs_ready (buffer116_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer117(
    .ins (buffer116_outs),
    .ins_valid (buffer116_outs_valid),
    .ins_ready (buffer116_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer117_outs),
    .outs_valid (buffer117_outs_valid),
    .outs_ready (buffer117_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork61(
    .ins (buffer117_outs),
    .ins_valid (buffer117_outs_valid),
    .ins_ready (buffer117_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork61_outs_1, fork61_outs_0}),
    .outs_valid ({fork61_outs_1_valid, fork61_outs_0_valid}),
    .outs_ready ({fork61_outs_1_ready, fork61_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi197(
    .ins (fork61_outs_0),
    .ins_valid (fork61_outs_0_valid),
    .ins_ready (fork61_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi197_outs),
    .outs_valid (extsi197_outs_valid),
    .outs_ready (extsi197_outs_ready)
  );

  oehb_dataless buffer118(
    .ins_valid (cond_br210_falseOut_valid),
    .ins_ready (cond_br210_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer118_outs_valid),
    .outs_ready (buffer118_outs_ready)
  );

  tehb_dataless buffer119(
    .ins_valid (buffer118_outs_valid),
    .ins_ready (buffer118_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer119_outs_valid),
    .outs_ready (buffer119_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork62(
    .ins_valid (buffer119_outs_valid),
    .ins_ready (buffer119_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork62_outs_6_valid, fork62_outs_5_valid, fork62_outs_4_valid, fork62_outs_3_valid, fork62_outs_2_valid, fork62_outs_1_valid, fork62_outs_0_valid}),
    .outs_ready ({fork62_outs_6_ready, fork62_outs_5_ready, fork62_outs_4_ready, fork62_outs_3_ready, fork62_outs_2_ready, fork62_outs_1_ready, fork62_outs_0_ready})
  );

  handshake_constant_140 #(.DATA_WIDTH(37)) constant363(
    .ctrl_valid (fork62_outs_5_valid),
    .ctrl_ready (fork62_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant363_outs),
    .outs_valid (constant363_outs_valid),
    .outs_ready (constant363_outs_ready)
  );

  handshake_constant_141 #(.DATA_WIDTH(29)) constant524(
    .ctrl_valid (fork62_outs_2_valid),
    .ctrl_ready (fork62_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant524_outs),
    .outs_valid (constant524_outs_valid),
    .outs_ready (constant524_outs_ready)
  );

  handshake_constant_142 #(.DATA_WIDTH(27)) constant365(
    .ctrl_valid (fork62_outs_4_valid),
    .ctrl_ready (fork62_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant365_outs),
    .outs_valid (constant365_outs_valid),
    .outs_ready (constant365_outs_ready)
  );

  handshake_constant_143 #(.DATA_WIDTH(20)) constant525(
    .ctrl_valid (fork62_outs_1_valid),
    .ctrl_ready (fork62_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant525_outs),
    .outs_valid (constant525_outs_valid),
    .outs_ready (constant525_outs_ready)
  );

  handshake_constant_144 #(.DATA_WIDTH(17)) constant367(
    .ctrl_valid (fork62_outs_3_valid),
    .ctrl_ready (fork62_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant367_outs),
    .outs_valid (constant367_outs_valid),
    .outs_ready (constant367_outs_ready)
  );

  handshake_constant_145 #(.DATA_WIDTH(7)) constant526(
    .ctrl_valid (fork62_outs_0_valid),
    .ctrl_ready (fork62_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant526_outs),
    .outs_valid (constant526_outs_valid),
    .outs_ready (constant526_outs_ready)
  );

  source source21(
    .clk (clk),
    .rst (rst),
    .outs_valid (source21_outs_valid),
    .outs_ready (source21_outs_ready)
  );

  handshake_constant_146 #(.DATA_WIDTH(6)) constant527(
    .ctrl_valid (source21_outs_valid),
    .ctrl_ready (source21_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant527_outs),
    .outs_valid (constant527_outs_valid),
    .outs_ready (constant527_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi20(
    .lhs (extsi197_outs),
    .lhs_valid (extsi197_outs_valid),
    .lhs_ready (extsi197_outs_ready),
    .rhs (constant527_outs),
    .rhs_valid (constant527_outs_valid),
    .rhs_ready (constant527_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi20_result),
    .result_valid (cmpi20_result_valid),
    .result_ready (cmpi20_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork63(
    .ins (cmpi20_result),
    .ins_valid (cmpi20_result_valid),
    .ins_ready (cmpi20_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork63_outs_8, fork63_outs_7, fork63_outs_6, fork63_outs_5, fork63_outs_4, fork63_outs_3, fork63_outs_2, fork63_outs_1, fork63_outs_0}),
    .outs_valid ({fork63_outs_8_valid, fork63_outs_7_valid, fork63_outs_6_valid, fork63_outs_5_valid, fork63_outs_4_valid, fork63_outs_3_valid, fork63_outs_2_valid, fork63_outs_1_valid, fork63_outs_0_valid}),
    .outs_ready ({fork63_outs_8_ready, fork63_outs_7_ready, fork63_outs_6_ready, fork63_outs_5_ready, fork63_outs_4_ready, fork63_outs_3_ready, fork63_outs_2_ready, fork63_outs_1_ready, fork63_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br212(
    .condition (fork63_outs_4),
    .condition_valid (fork63_outs_4_valid),
    .condition_ready (fork63_outs_4_ready),
    .data (constant363_outs),
    .data_valid (constant363_outs_valid),
    .data_ready (constant363_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br212_trueOut),
    .trueOut_valid (cond_br212_trueOut_valid),
    .trueOut_ready (cond_br212_trueOut_ready),
    .falseOut (cond_br212_falseOut),
    .falseOut_valid (cond_br212_falseOut_valid),
    .falseOut_ready (cond_br212_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink160(
    .ins (cond_br212_falseOut),
    .ins_valid (cond_br212_falseOut_valid),
    .ins_ready (cond_br212_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(29)) cond_br213(
    .condition (fork63_outs_7),
    .condition_valid (fork63_outs_7_valid),
    .condition_ready (fork63_outs_7_ready),
    .data (constant524_outs),
    .data_valid (constant524_outs_valid),
    .data_ready (constant524_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br213_trueOut),
    .trueOut_valid (cond_br213_trueOut_valid),
    .trueOut_ready (cond_br213_trueOut_ready),
    .falseOut (cond_br213_falseOut),
    .falseOut_valid (cond_br213_falseOut_valid),
    .falseOut_ready (cond_br213_falseOut_ready)
  );

  sink #(.DATA_TYPE(29)) sink161(
    .ins (cond_br213_falseOut),
    .ins_valid (cond_br213_falseOut_valid),
    .ins_ready (cond_br213_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(29), .OUTPUT_TYPE(33)) extsi198(
    .ins (cond_br213_trueOut),
    .ins_valid (cond_br213_trueOut_valid),
    .ins_ready (cond_br213_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi198_outs),
    .outs_valid (extsi198_outs_valid),
    .outs_ready (extsi198_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br214(
    .condition (fork63_outs_3),
    .condition_valid (fork63_outs_3_valid),
    .condition_ready (fork63_outs_3_ready),
    .data (constant365_outs),
    .data_valid (constant365_outs_valid),
    .data_ready (constant365_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br214_trueOut),
    .trueOut_valid (cond_br214_trueOut_valid),
    .trueOut_ready (cond_br214_trueOut_ready),
    .falseOut (cond_br214_falseOut),
    .falseOut_valid (cond_br214_falseOut_valid),
    .falseOut_ready (cond_br214_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink162(
    .ins (cond_br214_falseOut),
    .ins_valid (cond_br214_falseOut_valid),
    .ins_ready (cond_br214_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(20)) cond_br215(
    .condition (fork63_outs_6),
    .condition_valid (fork63_outs_6_valid),
    .condition_ready (fork63_outs_6_ready),
    .data (constant525_outs),
    .data_valid (constant525_outs_valid),
    .data_ready (constant525_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br215_trueOut),
    .trueOut_valid (cond_br215_trueOut_valid),
    .trueOut_ready (cond_br215_trueOut_ready),
    .falseOut (cond_br215_falseOut),
    .falseOut_valid (cond_br215_falseOut_valid),
    .falseOut_ready (cond_br215_falseOut_ready)
  );

  sink #(.DATA_TYPE(20)) sink163(
    .ins (cond_br215_falseOut),
    .ins_valid (cond_br215_falseOut_valid),
    .ins_ready (cond_br215_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(20), .OUTPUT_TYPE(22)) extsi199(
    .ins (cond_br215_trueOut),
    .ins_valid (cond_br215_trueOut_valid),
    .ins_ready (cond_br215_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi199_outs),
    .outs_valid (extsi199_outs_valid),
    .outs_ready (extsi199_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br216(
    .condition (fork63_outs_2),
    .condition_valid (fork63_outs_2_valid),
    .condition_ready (fork63_outs_2_ready),
    .data (constant367_outs),
    .data_valid (constant367_outs_valid),
    .data_ready (constant367_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br216_trueOut),
    .trueOut_valid (cond_br216_trueOut_valid),
    .trueOut_ready (cond_br216_trueOut_ready),
    .falseOut (cond_br216_falseOut),
    .falseOut_valid (cond_br216_falseOut_valid),
    .falseOut_ready (cond_br216_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink164(
    .ins (cond_br216_falseOut),
    .ins_valid (cond_br216_falseOut_valid),
    .ins_ready (cond_br216_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br217(
    .condition (fork63_outs_5),
    .condition_valid (fork63_outs_5_valid),
    .condition_ready (fork63_outs_5_ready),
    .data (constant526_outs),
    .data_valid (constant526_outs_valid),
    .data_ready (constant526_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br217_trueOut),
    .trueOut_valid (cond_br217_trueOut_valid),
    .trueOut_ready (cond_br217_trueOut_ready),
    .falseOut (cond_br217_falseOut),
    .falseOut_valid (cond_br217_falseOut_valid),
    .falseOut_ready (cond_br217_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink165(
    .ins (cond_br217_falseOut),
    .ins_valid (cond_br217_falseOut_valid),
    .ins_ready (cond_br217_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(12)) extsi200(
    .ins (cond_br217_trueOut),
    .ins_valid (cond_br217_trueOut_valid),
    .ins_ready (cond_br217_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi200_outs),
    .outs_valid (extsi200_outs_valid),
    .outs_ready (extsi200_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer114(
    .ins (cond_br209_falseOut),
    .ins_valid (cond_br209_falseOut_valid),
    .ins_ready (cond_br209_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer114_outs),
    .outs_valid (buffer114_outs_valid),
    .outs_ready (buffer114_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer115(
    .ins (buffer114_outs),
    .ins_valid (buffer114_outs_valid),
    .ins_ready (buffer114_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer115_outs),
    .outs_valid (buffer115_outs_valid),
    .outs_ready (buffer115_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br218(
    .condition (fork63_outs_0),
    .condition_valid (fork63_outs_0_valid),
    .condition_ready (fork63_outs_0_ready),
    .data (buffer115_outs),
    .data_valid (buffer115_outs_valid),
    .data_ready (buffer115_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br218_trueOut),
    .trueOut_valid (cond_br218_trueOut_valid),
    .trueOut_ready (cond_br218_trueOut_ready),
    .falseOut (cond_br218_falseOut),
    .falseOut_valid (cond_br218_falseOut_valid),
    .falseOut_ready (cond_br218_falseOut_ready)
  );

  cond_br_dataless cond_br219(
    .condition (fork63_outs_1),
    .condition_valid (fork63_outs_1_valid),
    .condition_ready (fork63_outs_1_ready),
    .data_valid (fork62_outs_6_valid),
    .data_ready (fork62_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br219_trueOut_valid),
    .trueOut_ready (cond_br219_trueOut_ready),
    .falseOut_valid (cond_br219_falseOut_valid),
    .falseOut_ready (cond_br219_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br220(
    .condition (fork63_outs_8),
    .condition_valid (fork63_outs_8_valid),
    .condition_ready (fork63_outs_8_ready),
    .data (fork61_outs_1),
    .data_valid (fork61_outs_1_valid),
    .data_ready (fork61_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br220_trueOut),
    .trueOut_valid (cond_br220_trueOut_valid),
    .trueOut_ready (cond_br220_trueOut_ready),
    .falseOut (cond_br220_falseOut),
    .falseOut_valid (cond_br220_falseOut_valid),
    .falseOut_ready (cond_br220_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink166(
    .ins (cond_br220_trueOut),
    .ins_valid (cond_br220_trueOut_valid),
    .ins_ready (cond_br220_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer122(
    .ins (cond_br220_falseOut),
    .ins_valid (cond_br220_falseOut_valid),
    .ins_ready (cond_br220_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer122_outs),
    .outs_valid (buffer122_outs_valid),
    .outs_ready (buffer122_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer123(
    .ins (buffer122_outs),
    .ins_valid (buffer122_outs_valid),
    .ins_ready (buffer122_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer123_outs),
    .outs_valid (buffer123_outs_valid),
    .outs_ready (buffer123_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork64(
    .ins (buffer123_outs),
    .ins_valid (buffer123_outs_valid),
    .ins_ready (buffer123_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork64_outs_1, fork64_outs_0}),
    .outs_valid ({fork64_outs_1_valid, fork64_outs_0_valid}),
    .outs_ready ({fork64_outs_1_ready, fork64_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi201(
    .ins (fork64_outs_0),
    .ins_valid (fork64_outs_0_valid),
    .ins_ready (fork64_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi201_outs),
    .outs_valid (extsi201_outs_valid),
    .outs_ready (extsi201_outs_ready)
  );

  oehb_dataless buffer124(
    .ins_valid (cond_br219_falseOut_valid),
    .ins_ready (cond_br219_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer124_outs_valid),
    .outs_ready (buffer124_outs_ready)
  );

  tehb_dataless buffer125(
    .ins_valid (buffer124_outs_valid),
    .ins_ready (buffer124_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer125_outs_valid),
    .outs_ready (buffer125_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork65(
    .ins_valid (buffer125_outs_valid),
    .ins_ready (buffer125_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork65_outs_6_valid, fork65_outs_5_valid, fork65_outs_4_valid, fork65_outs_3_valid, fork65_outs_2_valid, fork65_outs_1_valid, fork65_outs_0_valid}),
    .outs_ready ({fork65_outs_6_ready, fork65_outs_5_ready, fork65_outs_4_ready, fork65_outs_3_ready, fork65_outs_2_ready, fork65_outs_1_ready, fork65_outs_0_ready})
  );

  handshake_constant_147 #(.DATA_WIDTH(37)) constant370(
    .ctrl_valid (fork65_outs_5_valid),
    .ctrl_ready (fork65_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant370_outs),
    .outs_valid (constant370_outs_valid),
    .outs_ready (constant370_outs_ready)
  );

  handshake_constant_148 #(.DATA_WIDTH(29)) constant528(
    .ctrl_valid (fork65_outs_2_valid),
    .ctrl_ready (fork65_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant528_outs),
    .outs_valid (constant528_outs_valid),
    .outs_ready (constant528_outs_ready)
  );

  handshake_constant_149 #(.DATA_WIDTH(27)) constant372(
    .ctrl_valid (fork65_outs_4_valid),
    .ctrl_ready (fork65_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant372_outs),
    .outs_valid (constant372_outs_valid),
    .outs_ready (constant372_outs_ready)
  );

  handshake_constant_150 #(.DATA_WIDTH(19)) constant529(
    .ctrl_valid (fork65_outs_1_valid),
    .ctrl_ready (fork65_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant529_outs),
    .outs_valid (constant529_outs_valid),
    .outs_ready (constant529_outs_ready)
  );

  handshake_constant_151 #(.DATA_WIDTH(17)) constant374(
    .ctrl_valid (fork65_outs_3_valid),
    .ctrl_ready (fork65_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant374_outs),
    .outs_valid (constant374_outs_valid),
    .outs_ready (constant374_outs_ready)
  );

  handshake_constant_152 #(.DATA_WIDTH(8)) constant530(
    .ctrl_valid (fork65_outs_0_valid),
    .ctrl_ready (fork65_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant530_outs),
    .outs_valid (constant530_outs_valid),
    .outs_ready (constant530_outs_ready)
  );

  source source22(
    .clk (clk),
    .rst (rst),
    .outs_valid (source22_outs_valid),
    .outs_ready (source22_outs_ready)
  );

  handshake_constant_153 #(.DATA_WIDTH(6)) constant531(
    .ctrl_valid (source22_outs_valid),
    .ctrl_ready (source22_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant531_outs),
    .outs_valid (constant531_outs_valid),
    .outs_ready (constant531_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi21(
    .lhs (extsi201_outs),
    .lhs_valid (extsi201_outs_valid),
    .lhs_ready (extsi201_outs_ready),
    .rhs (constant531_outs),
    .rhs_valid (constant531_outs_valid),
    .rhs_ready (constant531_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi21_result),
    .result_valid (cmpi21_result_valid),
    .result_ready (cmpi21_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork66(
    .ins (cmpi21_result),
    .ins_valid (cmpi21_result_valid),
    .ins_ready (cmpi21_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork66_outs_8, fork66_outs_7, fork66_outs_6, fork66_outs_5, fork66_outs_4, fork66_outs_3, fork66_outs_2, fork66_outs_1, fork66_outs_0}),
    .outs_valid ({fork66_outs_8_valid, fork66_outs_7_valid, fork66_outs_6_valid, fork66_outs_5_valid, fork66_outs_4_valid, fork66_outs_3_valid, fork66_outs_2_valid, fork66_outs_1_valid, fork66_outs_0_valid}),
    .outs_ready ({fork66_outs_8_ready, fork66_outs_7_ready, fork66_outs_6_ready, fork66_outs_5_ready, fork66_outs_4_ready, fork66_outs_3_ready, fork66_outs_2_ready, fork66_outs_1_ready, fork66_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br221(
    .condition (fork66_outs_4),
    .condition_valid (fork66_outs_4_valid),
    .condition_ready (fork66_outs_4_ready),
    .data (constant370_outs),
    .data_valid (constant370_outs_valid),
    .data_ready (constant370_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br221_trueOut),
    .trueOut_valid (cond_br221_trueOut_valid),
    .trueOut_ready (cond_br221_trueOut_ready),
    .falseOut (cond_br221_falseOut),
    .falseOut_valid (cond_br221_falseOut_valid),
    .falseOut_ready (cond_br221_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink168(
    .ins (cond_br221_falseOut),
    .ins_valid (cond_br221_falseOut_valid),
    .ins_ready (cond_br221_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(29)) cond_br222(
    .condition (fork66_outs_7),
    .condition_valid (fork66_outs_7_valid),
    .condition_ready (fork66_outs_7_ready),
    .data (constant528_outs),
    .data_valid (constant528_outs_valid),
    .data_ready (constant528_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br222_trueOut),
    .trueOut_valid (cond_br222_trueOut_valid),
    .trueOut_ready (cond_br222_trueOut_ready),
    .falseOut (cond_br222_falseOut),
    .falseOut_valid (cond_br222_falseOut_valid),
    .falseOut_ready (cond_br222_falseOut_ready)
  );

  sink #(.DATA_TYPE(29)) sink169(
    .ins (cond_br222_falseOut),
    .ins_valid (cond_br222_falseOut_valid),
    .ins_ready (cond_br222_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(29), .OUTPUT_TYPE(33)) extsi202(
    .ins (cond_br222_trueOut),
    .ins_valid (cond_br222_trueOut_valid),
    .ins_ready (cond_br222_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi202_outs),
    .outs_valid (extsi202_outs_valid),
    .outs_ready (extsi202_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br223(
    .condition (fork66_outs_3),
    .condition_valid (fork66_outs_3_valid),
    .condition_ready (fork66_outs_3_ready),
    .data (constant372_outs),
    .data_valid (constant372_outs_valid),
    .data_ready (constant372_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br223_trueOut),
    .trueOut_valid (cond_br223_trueOut_valid),
    .trueOut_ready (cond_br223_trueOut_ready),
    .falseOut (cond_br223_falseOut),
    .falseOut_valid (cond_br223_falseOut_valid),
    .falseOut_ready (cond_br223_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink170(
    .ins (cond_br223_falseOut),
    .ins_valid (cond_br223_falseOut_valid),
    .ins_ready (cond_br223_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(19)) cond_br224(
    .condition (fork66_outs_6),
    .condition_valid (fork66_outs_6_valid),
    .condition_ready (fork66_outs_6_ready),
    .data (constant529_outs),
    .data_valid (constant529_outs_valid),
    .data_ready (constant529_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br224_trueOut),
    .trueOut_valid (cond_br224_trueOut_valid),
    .trueOut_ready (cond_br224_trueOut_ready),
    .falseOut (cond_br224_falseOut),
    .falseOut_valid (cond_br224_falseOut_valid),
    .falseOut_ready (cond_br224_falseOut_ready)
  );

  sink #(.DATA_TYPE(19)) sink171(
    .ins (cond_br224_falseOut),
    .ins_valid (cond_br224_falseOut_valid),
    .ins_ready (cond_br224_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(19), .OUTPUT_TYPE(22)) extsi203(
    .ins (cond_br224_trueOut),
    .ins_valid (cond_br224_trueOut_valid),
    .ins_ready (cond_br224_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi203_outs),
    .outs_valid (extsi203_outs_valid),
    .outs_ready (extsi203_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br225(
    .condition (fork66_outs_2),
    .condition_valid (fork66_outs_2_valid),
    .condition_ready (fork66_outs_2_ready),
    .data (constant374_outs),
    .data_valid (constant374_outs_valid),
    .data_ready (constant374_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br225_trueOut),
    .trueOut_valid (cond_br225_trueOut_valid),
    .trueOut_ready (cond_br225_trueOut_ready),
    .falseOut (cond_br225_falseOut),
    .falseOut_valid (cond_br225_falseOut_valid),
    .falseOut_ready (cond_br225_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink172(
    .ins (cond_br225_falseOut),
    .ins_valid (cond_br225_falseOut_valid),
    .ins_ready (cond_br225_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(8)) cond_br226(
    .condition (fork66_outs_5),
    .condition_valid (fork66_outs_5_valid),
    .condition_ready (fork66_outs_5_ready),
    .data (constant530_outs),
    .data_valid (constant530_outs_valid),
    .data_ready (constant530_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br226_trueOut),
    .trueOut_valid (cond_br226_trueOut_valid),
    .trueOut_ready (cond_br226_trueOut_ready),
    .falseOut (cond_br226_falseOut),
    .falseOut_valid (cond_br226_falseOut_valid),
    .falseOut_ready (cond_br226_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink173(
    .ins (cond_br226_falseOut),
    .ins_valid (cond_br226_falseOut_valid),
    .ins_ready (cond_br226_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(12)) extsi204(
    .ins (cond_br226_trueOut),
    .ins_valid (cond_br226_trueOut_valid),
    .ins_ready (cond_br226_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi204_outs),
    .outs_valid (extsi204_outs_valid),
    .outs_ready (extsi204_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer120(
    .ins (cond_br218_falseOut),
    .ins_valid (cond_br218_falseOut_valid),
    .ins_ready (cond_br218_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer120_outs),
    .outs_valid (buffer120_outs_valid),
    .outs_ready (buffer120_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer121(
    .ins (buffer120_outs),
    .ins_valid (buffer120_outs_valid),
    .ins_ready (buffer120_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer121_outs),
    .outs_valid (buffer121_outs_valid),
    .outs_ready (buffer121_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br227(
    .condition (fork66_outs_0),
    .condition_valid (fork66_outs_0_valid),
    .condition_ready (fork66_outs_0_ready),
    .data (buffer121_outs),
    .data_valid (buffer121_outs_valid),
    .data_ready (buffer121_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br227_trueOut),
    .trueOut_valid (cond_br227_trueOut_valid),
    .trueOut_ready (cond_br227_trueOut_ready),
    .falseOut (cond_br227_falseOut),
    .falseOut_valid (cond_br227_falseOut_valid),
    .falseOut_ready (cond_br227_falseOut_ready)
  );

  cond_br_dataless cond_br228(
    .condition (fork66_outs_1),
    .condition_valid (fork66_outs_1_valid),
    .condition_ready (fork66_outs_1_ready),
    .data_valid (fork65_outs_6_valid),
    .data_ready (fork65_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br228_trueOut_valid),
    .trueOut_ready (cond_br228_trueOut_ready),
    .falseOut_valid (cond_br228_falseOut_valid),
    .falseOut_ready (cond_br228_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br229(
    .condition (fork66_outs_8),
    .condition_valid (fork66_outs_8_valid),
    .condition_ready (fork66_outs_8_ready),
    .data (fork64_outs_1),
    .data_valid (fork64_outs_1_valid),
    .data_ready (fork64_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br229_trueOut),
    .trueOut_valid (cond_br229_trueOut_valid),
    .trueOut_ready (cond_br229_trueOut_ready),
    .falseOut (cond_br229_falseOut),
    .falseOut_valid (cond_br229_falseOut_valid),
    .falseOut_ready (cond_br229_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink174(
    .ins (cond_br229_trueOut),
    .ins_valid (cond_br229_trueOut_valid),
    .ins_ready (cond_br229_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer128(
    .ins (cond_br229_falseOut),
    .ins_valid (cond_br229_falseOut_valid),
    .ins_ready (cond_br229_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer128_outs),
    .outs_valid (buffer128_outs_valid),
    .outs_ready (buffer128_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer129(
    .ins (buffer128_outs),
    .ins_valid (buffer128_outs_valid),
    .ins_ready (buffer128_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer129_outs),
    .outs_valid (buffer129_outs_valid),
    .outs_ready (buffer129_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork67(
    .ins (buffer129_outs),
    .ins_valid (buffer129_outs_valid),
    .ins_ready (buffer129_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork67_outs_1, fork67_outs_0}),
    .outs_valid ({fork67_outs_1_valid, fork67_outs_0_valid}),
    .outs_ready ({fork67_outs_1_ready, fork67_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi205(
    .ins (fork67_outs_0),
    .ins_valid (fork67_outs_0_valid),
    .ins_ready (fork67_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi205_outs),
    .outs_valid (extsi205_outs_valid),
    .outs_ready (extsi205_outs_ready)
  );

  oehb_dataless buffer130(
    .ins_valid (cond_br228_falseOut_valid),
    .ins_ready (cond_br228_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer130_outs_valid),
    .outs_ready (buffer130_outs_ready)
  );

  tehb_dataless buffer131(
    .ins_valid (buffer130_outs_valid),
    .ins_ready (buffer130_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer131_outs_valid),
    .outs_ready (buffer131_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork68(
    .ins_valid (buffer131_outs_valid),
    .ins_ready (buffer131_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork68_outs_6_valid, fork68_outs_5_valid, fork68_outs_4_valid, fork68_outs_3_valid, fork68_outs_2_valid, fork68_outs_1_valid, fork68_outs_0_valid}),
    .outs_ready ({fork68_outs_6_ready, fork68_outs_5_ready, fork68_outs_4_ready, fork68_outs_3_ready, fork68_outs_2_ready, fork68_outs_1_ready, fork68_outs_0_ready})
  );

  handshake_constant_154 #(.DATA_WIDTH(37)) constant377(
    .ctrl_valid (fork68_outs_5_valid),
    .ctrl_ready (fork68_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant377_outs),
    .outs_valid (constant377_outs_valid),
    .outs_ready (constant377_outs_ready)
  );

  handshake_constant_155 #(.DATA_WIDTH(29)) constant532(
    .ctrl_valid (fork68_outs_2_valid),
    .ctrl_ready (fork68_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant532_outs),
    .outs_valid (constant532_outs_valid),
    .outs_ready (constant532_outs_ready)
  );

  handshake_constant_156 #(.DATA_WIDTH(27)) constant379(
    .ctrl_valid (fork68_outs_4_valid),
    .ctrl_ready (fork68_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant379_outs),
    .outs_valid (constant379_outs_valid),
    .outs_ready (constant379_outs_ready)
  );

  handshake_constant_157 #(.DATA_WIDTH(19)) constant533(
    .ctrl_valid (fork68_outs_1_valid),
    .ctrl_ready (fork68_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant533_outs),
    .outs_valid (constant533_outs_valid),
    .outs_ready (constant533_outs_ready)
  );

  handshake_constant_158 #(.DATA_WIDTH(17)) constant381(
    .ctrl_valid (fork68_outs_3_valid),
    .ctrl_ready (fork68_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant381_outs),
    .outs_valid (constant381_outs_valid),
    .outs_ready (constant381_outs_ready)
  );

  handshake_constant_159 #(.DATA_WIDTH(7)) constant534(
    .ctrl_valid (fork68_outs_0_valid),
    .ctrl_ready (fork68_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant534_outs),
    .outs_valid (constant534_outs_valid),
    .outs_ready (constant534_outs_ready)
  );

  source source23(
    .clk (clk),
    .rst (rst),
    .outs_valid (source23_outs_valid),
    .outs_ready (source23_outs_ready)
  );

  handshake_constant_160 #(.DATA_WIDTH(6)) constant535(
    .ctrl_valid (source23_outs_valid),
    .ctrl_ready (source23_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant535_outs),
    .outs_valid (constant535_outs_valid),
    .outs_ready (constant535_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi22(
    .lhs (extsi205_outs),
    .lhs_valid (extsi205_outs_valid),
    .lhs_ready (extsi205_outs_ready),
    .rhs (constant535_outs),
    .rhs_valid (constant535_outs_valid),
    .rhs_ready (constant535_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi22_result),
    .result_valid (cmpi22_result_valid),
    .result_ready (cmpi22_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork69(
    .ins (cmpi22_result),
    .ins_valid (cmpi22_result_valid),
    .ins_ready (cmpi22_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork69_outs_8, fork69_outs_7, fork69_outs_6, fork69_outs_5, fork69_outs_4, fork69_outs_3, fork69_outs_2, fork69_outs_1, fork69_outs_0}),
    .outs_valid ({fork69_outs_8_valid, fork69_outs_7_valid, fork69_outs_6_valid, fork69_outs_5_valid, fork69_outs_4_valid, fork69_outs_3_valid, fork69_outs_2_valid, fork69_outs_1_valid, fork69_outs_0_valid}),
    .outs_ready ({fork69_outs_8_ready, fork69_outs_7_ready, fork69_outs_6_ready, fork69_outs_5_ready, fork69_outs_4_ready, fork69_outs_3_ready, fork69_outs_2_ready, fork69_outs_1_ready, fork69_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br230(
    .condition (fork69_outs_4),
    .condition_valid (fork69_outs_4_valid),
    .condition_ready (fork69_outs_4_ready),
    .data (constant377_outs),
    .data_valid (constant377_outs_valid),
    .data_ready (constant377_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br230_trueOut),
    .trueOut_valid (cond_br230_trueOut_valid),
    .trueOut_ready (cond_br230_trueOut_ready),
    .falseOut (cond_br230_falseOut),
    .falseOut_valid (cond_br230_falseOut_valid),
    .falseOut_ready (cond_br230_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink176(
    .ins (cond_br230_falseOut),
    .ins_valid (cond_br230_falseOut_valid),
    .ins_ready (cond_br230_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(29)) cond_br231(
    .condition (fork69_outs_7),
    .condition_valid (fork69_outs_7_valid),
    .condition_ready (fork69_outs_7_ready),
    .data (constant532_outs),
    .data_valid (constant532_outs_valid),
    .data_ready (constant532_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br231_trueOut),
    .trueOut_valid (cond_br231_trueOut_valid),
    .trueOut_ready (cond_br231_trueOut_ready),
    .falseOut (cond_br231_falseOut),
    .falseOut_valid (cond_br231_falseOut_valid),
    .falseOut_ready (cond_br231_falseOut_ready)
  );

  sink #(.DATA_TYPE(29)) sink177(
    .ins (cond_br231_falseOut),
    .ins_valid (cond_br231_falseOut_valid),
    .ins_ready (cond_br231_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(29), .OUTPUT_TYPE(33)) extsi206(
    .ins (cond_br231_trueOut),
    .ins_valid (cond_br231_trueOut_valid),
    .ins_ready (cond_br231_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi206_outs),
    .outs_valid (extsi206_outs_valid),
    .outs_ready (extsi206_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br232(
    .condition (fork69_outs_3),
    .condition_valid (fork69_outs_3_valid),
    .condition_ready (fork69_outs_3_ready),
    .data (constant379_outs),
    .data_valid (constant379_outs_valid),
    .data_ready (constant379_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br232_trueOut),
    .trueOut_valid (cond_br232_trueOut_valid),
    .trueOut_ready (cond_br232_trueOut_ready),
    .falseOut (cond_br232_falseOut),
    .falseOut_valid (cond_br232_falseOut_valid),
    .falseOut_ready (cond_br232_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink178(
    .ins (cond_br232_falseOut),
    .ins_valid (cond_br232_falseOut_valid),
    .ins_ready (cond_br232_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(19)) cond_br233(
    .condition (fork69_outs_6),
    .condition_valid (fork69_outs_6_valid),
    .condition_ready (fork69_outs_6_ready),
    .data (constant533_outs),
    .data_valid (constant533_outs_valid),
    .data_ready (constant533_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br233_trueOut),
    .trueOut_valid (cond_br233_trueOut_valid),
    .trueOut_ready (cond_br233_trueOut_ready),
    .falseOut (cond_br233_falseOut),
    .falseOut_valid (cond_br233_falseOut_valid),
    .falseOut_ready (cond_br233_falseOut_ready)
  );

  sink #(.DATA_TYPE(19)) sink179(
    .ins (cond_br233_falseOut),
    .ins_valid (cond_br233_falseOut_valid),
    .ins_ready (cond_br233_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(19), .OUTPUT_TYPE(22)) extsi207(
    .ins (cond_br233_trueOut),
    .ins_valid (cond_br233_trueOut_valid),
    .ins_ready (cond_br233_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi207_outs),
    .outs_valid (extsi207_outs_valid),
    .outs_ready (extsi207_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br234(
    .condition (fork69_outs_2),
    .condition_valid (fork69_outs_2_valid),
    .condition_ready (fork69_outs_2_ready),
    .data (constant381_outs),
    .data_valid (constant381_outs_valid),
    .data_ready (constant381_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br234_trueOut),
    .trueOut_valid (cond_br234_trueOut_valid),
    .trueOut_ready (cond_br234_trueOut_ready),
    .falseOut (cond_br234_falseOut),
    .falseOut_valid (cond_br234_falseOut_valid),
    .falseOut_ready (cond_br234_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink180(
    .ins (cond_br234_falseOut),
    .ins_valid (cond_br234_falseOut_valid),
    .ins_ready (cond_br234_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br235(
    .condition (fork69_outs_5),
    .condition_valid (fork69_outs_5_valid),
    .condition_ready (fork69_outs_5_ready),
    .data (constant534_outs),
    .data_valid (constant534_outs_valid),
    .data_ready (constant534_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br235_trueOut),
    .trueOut_valid (cond_br235_trueOut_valid),
    .trueOut_ready (cond_br235_trueOut_ready),
    .falseOut (cond_br235_falseOut),
    .falseOut_valid (cond_br235_falseOut_valid),
    .falseOut_ready (cond_br235_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink181(
    .ins (cond_br235_falseOut),
    .ins_valid (cond_br235_falseOut_valid),
    .ins_ready (cond_br235_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(12)) extsi208(
    .ins (cond_br235_trueOut),
    .ins_valid (cond_br235_trueOut_valid),
    .ins_ready (cond_br235_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi208_outs),
    .outs_valid (extsi208_outs_valid),
    .outs_ready (extsi208_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer126(
    .ins (cond_br227_falseOut),
    .ins_valid (cond_br227_falseOut_valid),
    .ins_ready (cond_br227_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer126_outs),
    .outs_valid (buffer126_outs_valid),
    .outs_ready (buffer126_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer127(
    .ins (buffer126_outs),
    .ins_valid (buffer126_outs_valid),
    .ins_ready (buffer126_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer127_outs),
    .outs_valid (buffer127_outs_valid),
    .outs_ready (buffer127_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br236(
    .condition (fork69_outs_0),
    .condition_valid (fork69_outs_0_valid),
    .condition_ready (fork69_outs_0_ready),
    .data (buffer127_outs),
    .data_valid (buffer127_outs_valid),
    .data_ready (buffer127_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br236_trueOut),
    .trueOut_valid (cond_br236_trueOut_valid),
    .trueOut_ready (cond_br236_trueOut_ready),
    .falseOut (cond_br236_falseOut),
    .falseOut_valid (cond_br236_falseOut_valid),
    .falseOut_ready (cond_br236_falseOut_ready)
  );

  cond_br_dataless cond_br237(
    .condition (fork69_outs_1),
    .condition_valid (fork69_outs_1_valid),
    .condition_ready (fork69_outs_1_ready),
    .data_valid (fork68_outs_6_valid),
    .data_ready (fork68_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br237_trueOut_valid),
    .trueOut_ready (cond_br237_trueOut_ready),
    .falseOut_valid (cond_br237_falseOut_valid),
    .falseOut_ready (cond_br237_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br238(
    .condition (fork69_outs_8),
    .condition_valid (fork69_outs_8_valid),
    .condition_ready (fork69_outs_8_ready),
    .data (fork67_outs_1),
    .data_valid (fork67_outs_1_valid),
    .data_ready (fork67_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br238_trueOut),
    .trueOut_valid (cond_br238_trueOut_valid),
    .trueOut_ready (cond_br238_trueOut_ready),
    .falseOut (cond_br238_falseOut),
    .falseOut_valid (cond_br238_falseOut_valid),
    .falseOut_ready (cond_br238_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink182(
    .ins (cond_br238_trueOut),
    .ins_valid (cond_br238_trueOut_valid),
    .ins_ready (cond_br238_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer134(
    .ins (cond_br238_falseOut),
    .ins_valid (cond_br238_falseOut_valid),
    .ins_ready (cond_br238_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer134_outs),
    .outs_valid (buffer134_outs_valid),
    .outs_ready (buffer134_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer135(
    .ins (buffer134_outs),
    .ins_valid (buffer134_outs_valid),
    .ins_ready (buffer134_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer135_outs),
    .outs_valid (buffer135_outs_valid),
    .outs_ready (buffer135_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork70(
    .ins (buffer135_outs),
    .ins_valid (buffer135_outs_valid),
    .ins_ready (buffer135_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork70_outs_1, fork70_outs_0}),
    .outs_valid ({fork70_outs_1_valid, fork70_outs_0_valid}),
    .outs_ready ({fork70_outs_1_ready, fork70_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi209(
    .ins (fork70_outs_0),
    .ins_valid (fork70_outs_0_valid),
    .ins_ready (fork70_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi209_outs),
    .outs_valid (extsi209_outs_valid),
    .outs_ready (extsi209_outs_ready)
  );

  oehb_dataless buffer136(
    .ins_valid (cond_br237_falseOut_valid),
    .ins_ready (cond_br237_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer136_outs_valid),
    .outs_ready (buffer136_outs_ready)
  );

  tehb_dataless buffer137(
    .ins_valid (buffer136_outs_valid),
    .ins_ready (buffer136_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer137_outs_valid),
    .outs_ready (buffer137_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork71(
    .ins_valid (buffer137_outs_valid),
    .ins_ready (buffer137_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork71_outs_6_valid, fork71_outs_5_valid, fork71_outs_4_valid, fork71_outs_3_valid, fork71_outs_2_valid, fork71_outs_1_valid, fork71_outs_0_valid}),
    .outs_ready ({fork71_outs_6_ready, fork71_outs_5_ready, fork71_outs_4_ready, fork71_outs_3_ready, fork71_outs_2_ready, fork71_outs_1_ready, fork71_outs_0_ready})
  );

  handshake_constant_138 #(.DATA_WIDTH(7)) constant536(
    .ctrl_valid (fork71_outs_2_valid),
    .ctrl_ready (fork71_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant536_outs),
    .outs_valid (constant536_outs_valid),
    .outs_ready (constant536_outs_ready)
  );

  handshake_constant_161 #(.DATA_WIDTH(37)) constant385(
    .ctrl_valid (fork71_outs_5_valid),
    .ctrl_ready (fork71_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant385_outs),
    .outs_valid (constant385_outs_valid),
    .outs_ready (constant385_outs_ready)
  );

  handshake_constant_162 #(.DATA_WIDTH(29)) constant537(
    .ctrl_valid (fork71_outs_1_valid),
    .ctrl_ready (fork71_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant537_outs),
    .outs_valid (constant537_outs_valid),
    .outs_ready (constant537_outs_ready)
  );

  handshake_constant_163 #(.DATA_WIDTH(27)) constant387(
    .ctrl_valid (fork71_outs_4_valid),
    .ctrl_ready (fork71_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant387_outs),
    .outs_valid (constant387_outs_valid),
    .outs_ready (constant387_outs_ready)
  );

  handshake_constant_164 #(.DATA_WIDTH(19)) constant538(
    .ctrl_valid (fork71_outs_0_valid),
    .ctrl_ready (fork71_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant538_outs),
    .outs_valid (constant538_outs_valid),
    .outs_ready (constant538_outs_ready)
  );

  handshake_constant_165 #(.DATA_WIDTH(17)) constant389(
    .ctrl_valid (fork71_outs_3_valid),
    .ctrl_ready (fork71_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant389_outs),
    .outs_valid (constant389_outs_valid),
    .outs_ready (constant389_outs_ready)
  );

  source source24(
    .clk (clk),
    .rst (rst),
    .outs_valid (source24_outs_valid),
    .outs_ready (source24_outs_ready)
  );

  handshake_constant_166 #(.DATA_WIDTH(6)) constant539(
    .ctrl_valid (source24_outs_valid),
    .ctrl_ready (source24_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant539_outs),
    .outs_valid (constant539_outs_valid),
    .outs_ready (constant539_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi23(
    .lhs (extsi209_outs),
    .lhs_valid (extsi209_outs_valid),
    .lhs_ready (extsi209_outs_ready),
    .rhs (constant539_outs),
    .rhs_valid (constant539_outs_valid),
    .rhs_ready (constant539_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi23_result),
    .result_valid (cmpi23_result_valid),
    .result_ready (cmpi23_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork72(
    .ins (cmpi23_result),
    .ins_valid (cmpi23_result_valid),
    .ins_ready (cmpi23_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork72_outs_8, fork72_outs_7, fork72_outs_6, fork72_outs_5, fork72_outs_4, fork72_outs_3, fork72_outs_2, fork72_outs_1, fork72_outs_0}),
    .outs_valid ({fork72_outs_8_valid, fork72_outs_7_valid, fork72_outs_6_valid, fork72_outs_5_valid, fork72_outs_4_valid, fork72_outs_3_valid, fork72_outs_2_valid, fork72_outs_1_valid, fork72_outs_0_valid}),
    .outs_ready ({fork72_outs_8_ready, fork72_outs_7_ready, fork72_outs_6_ready, fork72_outs_5_ready, fork72_outs_4_ready, fork72_outs_3_ready, fork72_outs_2_ready, fork72_outs_1_ready, fork72_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br239(
    .condition (fork72_outs_4),
    .condition_valid (fork72_outs_4_valid),
    .condition_ready (fork72_outs_4_ready),
    .data (constant385_outs),
    .data_valid (constant385_outs_valid),
    .data_ready (constant385_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br239_trueOut),
    .trueOut_valid (cond_br239_trueOut_valid),
    .trueOut_ready (cond_br239_trueOut_ready),
    .falseOut (cond_br239_falseOut),
    .falseOut_valid (cond_br239_falseOut_valid),
    .falseOut_ready (cond_br239_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink184(
    .ins (cond_br239_falseOut),
    .ins_valid (cond_br239_falseOut_valid),
    .ins_ready (cond_br239_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(29)) cond_br240(
    .condition (fork72_outs_7),
    .condition_valid (fork72_outs_7_valid),
    .condition_ready (fork72_outs_7_ready),
    .data (constant537_outs),
    .data_valid (constant537_outs_valid),
    .data_ready (constant537_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br240_trueOut),
    .trueOut_valid (cond_br240_trueOut_valid),
    .trueOut_ready (cond_br240_trueOut_ready),
    .falseOut (cond_br240_falseOut),
    .falseOut_valid (cond_br240_falseOut_valid),
    .falseOut_ready (cond_br240_falseOut_ready)
  );

  sink #(.DATA_TYPE(29)) sink185(
    .ins (cond_br240_falseOut),
    .ins_valid (cond_br240_falseOut_valid),
    .ins_ready (cond_br240_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(29), .OUTPUT_TYPE(33)) extsi210(
    .ins (cond_br240_trueOut),
    .ins_valid (cond_br240_trueOut_valid),
    .ins_ready (cond_br240_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi210_outs),
    .outs_valid (extsi210_outs_valid),
    .outs_ready (extsi210_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br241(
    .condition (fork72_outs_3),
    .condition_valid (fork72_outs_3_valid),
    .condition_ready (fork72_outs_3_ready),
    .data (constant387_outs),
    .data_valid (constant387_outs_valid),
    .data_ready (constant387_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br241_trueOut),
    .trueOut_valid (cond_br241_trueOut_valid),
    .trueOut_ready (cond_br241_trueOut_ready),
    .falseOut (cond_br241_falseOut),
    .falseOut_valid (cond_br241_falseOut_valid),
    .falseOut_ready (cond_br241_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink186(
    .ins (cond_br241_falseOut),
    .ins_valid (cond_br241_falseOut_valid),
    .ins_ready (cond_br241_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(19)) cond_br242(
    .condition (fork72_outs_6),
    .condition_valid (fork72_outs_6_valid),
    .condition_ready (fork72_outs_6_ready),
    .data (constant538_outs),
    .data_valid (constant538_outs_valid),
    .data_ready (constant538_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br242_trueOut),
    .trueOut_valid (cond_br242_trueOut_valid),
    .trueOut_ready (cond_br242_trueOut_ready),
    .falseOut (cond_br242_falseOut),
    .falseOut_valid (cond_br242_falseOut_valid),
    .falseOut_ready (cond_br242_falseOut_ready)
  );

  sink #(.DATA_TYPE(19)) sink187(
    .ins (cond_br242_falseOut),
    .ins_valid (cond_br242_falseOut_valid),
    .ins_ready (cond_br242_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(19), .OUTPUT_TYPE(22)) extsi211(
    .ins (cond_br242_trueOut),
    .ins_valid (cond_br242_trueOut_valid),
    .ins_ready (cond_br242_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi211_outs),
    .outs_valid (extsi211_outs_valid),
    .outs_ready (extsi211_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br243(
    .condition (fork72_outs_2),
    .condition_valid (fork72_outs_2_valid),
    .condition_ready (fork72_outs_2_ready),
    .data (constant389_outs),
    .data_valid (constant389_outs_valid),
    .data_ready (constant389_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br243_trueOut),
    .trueOut_valid (cond_br243_trueOut_valid),
    .trueOut_ready (cond_br243_trueOut_ready),
    .falseOut (cond_br243_falseOut),
    .falseOut_valid (cond_br243_falseOut_valid),
    .falseOut_ready (cond_br243_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink188(
    .ins (cond_br243_falseOut),
    .ins_valid (cond_br243_falseOut_valid),
    .ins_ready (cond_br243_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br244(
    .condition (fork72_outs_5),
    .condition_valid (fork72_outs_5_valid),
    .condition_ready (fork72_outs_5_ready),
    .data (constant536_outs),
    .data_valid (constant536_outs_valid),
    .data_ready (constant536_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br244_trueOut),
    .trueOut_valid (cond_br244_trueOut_valid),
    .trueOut_ready (cond_br244_trueOut_ready),
    .falseOut (cond_br244_falseOut),
    .falseOut_valid (cond_br244_falseOut_valid),
    .falseOut_ready (cond_br244_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink189(
    .ins (cond_br244_falseOut),
    .ins_valid (cond_br244_falseOut_valid),
    .ins_ready (cond_br244_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(12)) extsi212(
    .ins (cond_br244_trueOut),
    .ins_valid (cond_br244_trueOut_valid),
    .ins_ready (cond_br244_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi212_outs),
    .outs_valid (extsi212_outs_valid),
    .outs_ready (extsi212_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer132(
    .ins (cond_br236_falseOut),
    .ins_valid (cond_br236_falseOut_valid),
    .ins_ready (cond_br236_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer132_outs),
    .outs_valid (buffer132_outs_valid),
    .outs_ready (buffer132_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer133(
    .ins (buffer132_outs),
    .ins_valid (buffer132_outs_valid),
    .ins_ready (buffer132_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer133_outs),
    .outs_valid (buffer133_outs_valid),
    .outs_ready (buffer133_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br245(
    .condition (fork72_outs_0),
    .condition_valid (fork72_outs_0_valid),
    .condition_ready (fork72_outs_0_ready),
    .data (buffer133_outs),
    .data_valid (buffer133_outs_valid),
    .data_ready (buffer133_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br245_trueOut),
    .trueOut_valid (cond_br245_trueOut_valid),
    .trueOut_ready (cond_br245_trueOut_ready),
    .falseOut (cond_br245_falseOut),
    .falseOut_valid (cond_br245_falseOut_valid),
    .falseOut_ready (cond_br245_falseOut_ready)
  );

  cond_br_dataless cond_br246(
    .condition (fork72_outs_1),
    .condition_valid (fork72_outs_1_valid),
    .condition_ready (fork72_outs_1_ready),
    .data_valid (fork71_outs_6_valid),
    .data_ready (fork71_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br246_trueOut_valid),
    .trueOut_ready (cond_br246_trueOut_ready),
    .falseOut_valid (cond_br246_falseOut_valid),
    .falseOut_ready (cond_br246_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br247(
    .condition (fork72_outs_8),
    .condition_valid (fork72_outs_8_valid),
    .condition_ready (fork72_outs_8_ready),
    .data (fork70_outs_1),
    .data_valid (fork70_outs_1_valid),
    .data_ready (fork70_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br247_trueOut),
    .trueOut_valid (cond_br247_trueOut_valid),
    .trueOut_ready (cond_br247_trueOut_ready),
    .falseOut (cond_br247_falseOut),
    .falseOut_valid (cond_br247_falseOut_valid),
    .falseOut_ready (cond_br247_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink190(
    .ins (cond_br247_trueOut),
    .ins_valid (cond_br247_trueOut_valid),
    .ins_ready (cond_br247_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer140(
    .ins (cond_br247_falseOut),
    .ins_valid (cond_br247_falseOut_valid),
    .ins_ready (cond_br247_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer140_outs),
    .outs_valid (buffer140_outs_valid),
    .outs_ready (buffer140_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer141(
    .ins (buffer140_outs),
    .ins_valid (buffer140_outs_valid),
    .ins_ready (buffer140_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer141_outs),
    .outs_valid (buffer141_outs_valid),
    .outs_ready (buffer141_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork73(
    .ins (buffer141_outs),
    .ins_valid (buffer141_outs_valid),
    .ins_ready (buffer141_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork73_outs_1, fork73_outs_0}),
    .outs_valid ({fork73_outs_1_valid, fork73_outs_0_valid}),
    .outs_ready ({fork73_outs_1_ready, fork73_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi213(
    .ins (fork73_outs_0),
    .ins_valid (fork73_outs_0_valid),
    .ins_ready (fork73_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi213_outs),
    .outs_valid (extsi213_outs_valid),
    .outs_ready (extsi213_outs_ready)
  );

  oehb_dataless buffer142(
    .ins_valid (cond_br246_falseOut_valid),
    .ins_ready (cond_br246_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer142_outs_valid),
    .outs_ready (buffer142_outs_ready)
  );

  tehb_dataless buffer143(
    .ins_valid (buffer142_outs_valid),
    .ins_ready (buffer142_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer143_outs_valid),
    .outs_ready (buffer143_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork74(
    .ins_valid (buffer143_outs_valid),
    .ins_ready (buffer143_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork74_outs_6_valid, fork74_outs_5_valid, fork74_outs_4_valid, fork74_outs_3_valid, fork74_outs_2_valid, fork74_outs_1_valid, fork74_outs_0_valid}),
    .outs_ready ({fork74_outs_6_ready, fork74_outs_5_ready, fork74_outs_4_ready, fork74_outs_3_ready, fork74_outs_2_ready, fork74_outs_1_ready, fork74_outs_0_ready})
  );

  handshake_constant_167 #(.DATA_WIDTH(37)) constant391(
    .ctrl_valid (fork74_outs_5_valid),
    .ctrl_ready (fork74_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant391_outs),
    .outs_valid (constant391_outs_valid),
    .outs_ready (constant391_outs_ready)
  );

  handshake_constant_168 #(.DATA_WIDTH(28)) constant540(
    .ctrl_valid (fork74_outs_2_valid),
    .ctrl_ready (fork74_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant540_outs),
    .outs_valid (constant540_outs_valid),
    .outs_ready (constant540_outs_ready)
  );

  handshake_constant_169 #(.DATA_WIDTH(27)) constant393(
    .ctrl_valid (fork74_outs_4_valid),
    .ctrl_ready (fork74_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant393_outs),
    .outs_valid (constant393_outs_valid),
    .outs_ready (constant393_outs_ready)
  );

  handshake_constant_170 #(.DATA_WIDTH(19)) constant541(
    .ctrl_valid (fork74_outs_1_valid),
    .ctrl_ready (fork74_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant541_outs),
    .outs_valid (constant541_outs_valid),
    .outs_ready (constant541_outs_ready)
  );

  handshake_constant_171 #(.DATA_WIDTH(17)) constant395(
    .ctrl_valid (fork74_outs_3_valid),
    .ctrl_ready (fork74_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant395_outs),
    .outs_valid (constant395_outs_valid),
    .outs_ready (constant395_outs_ready)
  );

  handshake_constant_172 #(.DATA_WIDTH(7)) constant542(
    .ctrl_valid (fork74_outs_0_valid),
    .ctrl_ready (fork74_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant542_outs),
    .outs_valid (constant542_outs_valid),
    .outs_ready (constant542_outs_ready)
  );

  source source25(
    .clk (clk),
    .rst (rst),
    .outs_valid (source25_outs_valid),
    .outs_ready (source25_outs_ready)
  );

  handshake_constant_173 #(.DATA_WIDTH(6)) constant543(
    .ctrl_valid (source25_outs_valid),
    .ctrl_ready (source25_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant543_outs),
    .outs_valid (constant543_outs_valid),
    .outs_ready (constant543_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi24(
    .lhs (extsi213_outs),
    .lhs_valid (extsi213_outs_valid),
    .lhs_ready (extsi213_outs_ready),
    .rhs (constant543_outs),
    .rhs_valid (constant543_outs_valid),
    .rhs_ready (constant543_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi24_result),
    .result_valid (cmpi24_result_valid),
    .result_ready (cmpi24_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork75(
    .ins (cmpi24_result),
    .ins_valid (cmpi24_result_valid),
    .ins_ready (cmpi24_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork75_outs_8, fork75_outs_7, fork75_outs_6, fork75_outs_5, fork75_outs_4, fork75_outs_3, fork75_outs_2, fork75_outs_1, fork75_outs_0}),
    .outs_valid ({fork75_outs_8_valid, fork75_outs_7_valid, fork75_outs_6_valid, fork75_outs_5_valid, fork75_outs_4_valid, fork75_outs_3_valid, fork75_outs_2_valid, fork75_outs_1_valid, fork75_outs_0_valid}),
    .outs_ready ({fork75_outs_8_ready, fork75_outs_7_ready, fork75_outs_6_ready, fork75_outs_5_ready, fork75_outs_4_ready, fork75_outs_3_ready, fork75_outs_2_ready, fork75_outs_1_ready, fork75_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br248(
    .condition (fork75_outs_4),
    .condition_valid (fork75_outs_4_valid),
    .condition_ready (fork75_outs_4_ready),
    .data (constant391_outs),
    .data_valid (constant391_outs_valid),
    .data_ready (constant391_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br248_trueOut),
    .trueOut_valid (cond_br248_trueOut_valid),
    .trueOut_ready (cond_br248_trueOut_ready),
    .falseOut (cond_br248_falseOut),
    .falseOut_valid (cond_br248_falseOut_valid),
    .falseOut_ready (cond_br248_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink192(
    .ins (cond_br248_falseOut),
    .ins_valid (cond_br248_falseOut_valid),
    .ins_ready (cond_br248_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(28)) cond_br249(
    .condition (fork75_outs_7),
    .condition_valid (fork75_outs_7_valid),
    .condition_ready (fork75_outs_7_ready),
    .data (constant540_outs),
    .data_valid (constant540_outs_valid),
    .data_ready (constant540_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br249_trueOut),
    .trueOut_valid (cond_br249_trueOut_valid),
    .trueOut_ready (cond_br249_trueOut_ready),
    .falseOut (cond_br249_falseOut),
    .falseOut_valid (cond_br249_falseOut_valid),
    .falseOut_ready (cond_br249_falseOut_ready)
  );

  sink #(.DATA_TYPE(28)) sink193(
    .ins (cond_br249_falseOut),
    .ins_valid (cond_br249_falseOut_valid),
    .ins_ready (cond_br249_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(28), .OUTPUT_TYPE(33)) extsi214(
    .ins (cond_br249_trueOut),
    .ins_valid (cond_br249_trueOut_valid),
    .ins_ready (cond_br249_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi214_outs),
    .outs_valid (extsi214_outs_valid),
    .outs_ready (extsi214_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br250(
    .condition (fork75_outs_3),
    .condition_valid (fork75_outs_3_valid),
    .condition_ready (fork75_outs_3_ready),
    .data (constant393_outs),
    .data_valid (constant393_outs_valid),
    .data_ready (constant393_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br250_trueOut),
    .trueOut_valid (cond_br250_trueOut_valid),
    .trueOut_ready (cond_br250_trueOut_ready),
    .falseOut (cond_br250_falseOut),
    .falseOut_valid (cond_br250_falseOut_valid),
    .falseOut_ready (cond_br250_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink194(
    .ins (cond_br250_falseOut),
    .ins_valid (cond_br250_falseOut_valid),
    .ins_ready (cond_br250_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(19)) cond_br251(
    .condition (fork75_outs_6),
    .condition_valid (fork75_outs_6_valid),
    .condition_ready (fork75_outs_6_ready),
    .data (constant541_outs),
    .data_valid (constant541_outs_valid),
    .data_ready (constant541_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br251_trueOut),
    .trueOut_valid (cond_br251_trueOut_valid),
    .trueOut_ready (cond_br251_trueOut_ready),
    .falseOut (cond_br251_falseOut),
    .falseOut_valid (cond_br251_falseOut_valid),
    .falseOut_ready (cond_br251_falseOut_ready)
  );

  sink #(.DATA_TYPE(19)) sink195(
    .ins (cond_br251_falseOut),
    .ins_valid (cond_br251_falseOut_valid),
    .ins_ready (cond_br251_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(19), .OUTPUT_TYPE(22)) extsi215(
    .ins (cond_br251_trueOut),
    .ins_valid (cond_br251_trueOut_valid),
    .ins_ready (cond_br251_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi215_outs),
    .outs_valid (extsi215_outs_valid),
    .outs_ready (extsi215_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br252(
    .condition (fork75_outs_2),
    .condition_valid (fork75_outs_2_valid),
    .condition_ready (fork75_outs_2_ready),
    .data (constant395_outs),
    .data_valid (constant395_outs_valid),
    .data_ready (constant395_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br252_trueOut),
    .trueOut_valid (cond_br252_trueOut_valid),
    .trueOut_ready (cond_br252_trueOut_ready),
    .falseOut (cond_br252_falseOut),
    .falseOut_valid (cond_br252_falseOut_valid),
    .falseOut_ready (cond_br252_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink196(
    .ins (cond_br252_falseOut),
    .ins_valid (cond_br252_falseOut_valid),
    .ins_ready (cond_br252_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br253(
    .condition (fork75_outs_5),
    .condition_valid (fork75_outs_5_valid),
    .condition_ready (fork75_outs_5_ready),
    .data (constant542_outs),
    .data_valid (constant542_outs_valid),
    .data_ready (constant542_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br253_trueOut),
    .trueOut_valid (cond_br253_trueOut_valid),
    .trueOut_ready (cond_br253_trueOut_ready),
    .falseOut (cond_br253_falseOut),
    .falseOut_valid (cond_br253_falseOut_valid),
    .falseOut_ready (cond_br253_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink197(
    .ins (cond_br253_falseOut),
    .ins_valid (cond_br253_falseOut_valid),
    .ins_ready (cond_br253_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(12)) extsi216(
    .ins (cond_br253_trueOut),
    .ins_valid (cond_br253_trueOut_valid),
    .ins_ready (cond_br253_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi216_outs),
    .outs_valid (extsi216_outs_valid),
    .outs_ready (extsi216_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer138(
    .ins (cond_br245_falseOut),
    .ins_valid (cond_br245_falseOut_valid),
    .ins_ready (cond_br245_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer138_outs),
    .outs_valid (buffer138_outs_valid),
    .outs_ready (buffer138_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer139(
    .ins (buffer138_outs),
    .ins_valid (buffer138_outs_valid),
    .ins_ready (buffer138_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer139_outs),
    .outs_valid (buffer139_outs_valid),
    .outs_ready (buffer139_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br254(
    .condition (fork75_outs_0),
    .condition_valid (fork75_outs_0_valid),
    .condition_ready (fork75_outs_0_ready),
    .data (buffer139_outs),
    .data_valid (buffer139_outs_valid),
    .data_ready (buffer139_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br254_trueOut),
    .trueOut_valid (cond_br254_trueOut_valid),
    .trueOut_ready (cond_br254_trueOut_ready),
    .falseOut (cond_br254_falseOut),
    .falseOut_valid (cond_br254_falseOut_valid),
    .falseOut_ready (cond_br254_falseOut_ready)
  );

  cond_br_dataless cond_br255(
    .condition (fork75_outs_1),
    .condition_valid (fork75_outs_1_valid),
    .condition_ready (fork75_outs_1_ready),
    .data_valid (fork74_outs_6_valid),
    .data_ready (fork74_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br255_trueOut_valid),
    .trueOut_ready (cond_br255_trueOut_ready),
    .falseOut_valid (cond_br255_falseOut_valid),
    .falseOut_ready (cond_br255_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br256(
    .condition (fork75_outs_8),
    .condition_valid (fork75_outs_8_valid),
    .condition_ready (fork75_outs_8_ready),
    .data (fork73_outs_1),
    .data_valid (fork73_outs_1_valid),
    .data_ready (fork73_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br256_trueOut),
    .trueOut_valid (cond_br256_trueOut_valid),
    .trueOut_ready (cond_br256_trueOut_ready),
    .falseOut (cond_br256_falseOut),
    .falseOut_valid (cond_br256_falseOut_valid),
    .falseOut_ready (cond_br256_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink198(
    .ins (cond_br256_trueOut),
    .ins_valid (cond_br256_trueOut_valid),
    .ins_ready (cond_br256_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer146(
    .ins (cond_br256_falseOut),
    .ins_valid (cond_br256_falseOut_valid),
    .ins_ready (cond_br256_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer146_outs),
    .outs_valid (buffer146_outs_valid),
    .outs_ready (buffer146_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer147(
    .ins (buffer146_outs),
    .ins_valid (buffer146_outs_valid),
    .ins_ready (buffer146_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer147_outs),
    .outs_valid (buffer147_outs_valid),
    .outs_ready (buffer147_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork76(
    .ins (buffer147_outs),
    .ins_valid (buffer147_outs_valid),
    .ins_ready (buffer147_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork76_outs_1, fork76_outs_0}),
    .outs_valid ({fork76_outs_1_valid, fork76_outs_0_valid}),
    .outs_ready ({fork76_outs_1_ready, fork76_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi217(
    .ins (fork76_outs_0),
    .ins_valid (fork76_outs_0_valid),
    .ins_ready (fork76_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi217_outs),
    .outs_valid (extsi217_outs_valid),
    .outs_ready (extsi217_outs_ready)
  );

  oehb_dataless buffer148(
    .ins_valid (cond_br255_falseOut_valid),
    .ins_ready (cond_br255_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer148_outs_valid),
    .outs_ready (buffer148_outs_ready)
  );

  tehb_dataless buffer149(
    .ins_valid (buffer148_outs_valid),
    .ins_ready (buffer148_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer149_outs_valid),
    .outs_ready (buffer149_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork77(
    .ins_valid (buffer149_outs_valid),
    .ins_ready (buffer149_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork77_outs_6_valid, fork77_outs_5_valid, fork77_outs_4_valid, fork77_outs_3_valid, fork77_outs_2_valid, fork77_outs_1_valid, fork77_outs_0_valid}),
    .outs_ready ({fork77_outs_6_ready, fork77_outs_5_ready, fork77_outs_4_ready, fork77_outs_3_ready, fork77_outs_2_ready, fork77_outs_1_ready, fork77_outs_0_ready})
  );

  handshake_constant_174 #(.DATA_WIDTH(37)) constant398(
    .ctrl_valid (fork77_outs_5_valid),
    .ctrl_ready (fork77_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant398_outs),
    .outs_valid (constant398_outs_valid),
    .outs_ready (constant398_outs_ready)
  );

  handshake_constant_175 #(.DATA_WIDTH(28)) constant544(
    .ctrl_valid (fork77_outs_2_valid),
    .ctrl_ready (fork77_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant544_outs),
    .outs_valid (constant544_outs_valid),
    .outs_ready (constant544_outs_ready)
  );

  handshake_constant_176 #(.DATA_WIDTH(27)) constant400(
    .ctrl_valid (fork77_outs_4_valid),
    .ctrl_ready (fork77_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant400_outs),
    .outs_valid (constant400_outs_valid),
    .outs_ready (constant400_outs_ready)
  );

  handshake_constant_177 #(.DATA_WIDTH(18)) constant545(
    .ctrl_valid (fork77_outs_1_valid),
    .ctrl_ready (fork77_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant545_outs),
    .outs_valid (constant545_outs_valid),
    .outs_ready (constant545_outs_ready)
  );

  handshake_constant_178 #(.DATA_WIDTH(17)) constant402(
    .ctrl_valid (fork77_outs_3_valid),
    .ctrl_ready (fork77_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant402_outs),
    .outs_valid (constant402_outs_valid),
    .outs_ready (constant402_outs_ready)
  );

  handshake_constant_179 #(.DATA_WIDTH(7)) constant546(
    .ctrl_valid (fork77_outs_0_valid),
    .ctrl_ready (fork77_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant546_outs),
    .outs_valid (constant546_outs_valid),
    .outs_ready (constant546_outs_ready)
  );

  source source26(
    .clk (clk),
    .rst (rst),
    .outs_valid (source26_outs_valid),
    .outs_ready (source26_outs_ready)
  );

  handshake_constant_180 #(.DATA_WIDTH(6)) constant547(
    .ctrl_valid (source26_outs_valid),
    .ctrl_ready (source26_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant547_outs),
    .outs_valid (constant547_outs_valid),
    .outs_ready (constant547_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi25(
    .lhs (extsi217_outs),
    .lhs_valid (extsi217_outs_valid),
    .lhs_ready (extsi217_outs_ready),
    .rhs (constant547_outs),
    .rhs_valid (constant547_outs_valid),
    .rhs_ready (constant547_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi25_result),
    .result_valid (cmpi25_result_valid),
    .result_ready (cmpi25_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork78(
    .ins (cmpi25_result),
    .ins_valid (cmpi25_result_valid),
    .ins_ready (cmpi25_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork78_outs_8, fork78_outs_7, fork78_outs_6, fork78_outs_5, fork78_outs_4, fork78_outs_3, fork78_outs_2, fork78_outs_1, fork78_outs_0}),
    .outs_valid ({fork78_outs_8_valid, fork78_outs_7_valid, fork78_outs_6_valid, fork78_outs_5_valid, fork78_outs_4_valid, fork78_outs_3_valid, fork78_outs_2_valid, fork78_outs_1_valid, fork78_outs_0_valid}),
    .outs_ready ({fork78_outs_8_ready, fork78_outs_7_ready, fork78_outs_6_ready, fork78_outs_5_ready, fork78_outs_4_ready, fork78_outs_3_ready, fork78_outs_2_ready, fork78_outs_1_ready, fork78_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br257(
    .condition (fork78_outs_4),
    .condition_valid (fork78_outs_4_valid),
    .condition_ready (fork78_outs_4_ready),
    .data (constant398_outs),
    .data_valid (constant398_outs_valid),
    .data_ready (constant398_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br257_trueOut),
    .trueOut_valid (cond_br257_trueOut_valid),
    .trueOut_ready (cond_br257_trueOut_ready),
    .falseOut (cond_br257_falseOut),
    .falseOut_valid (cond_br257_falseOut_valid),
    .falseOut_ready (cond_br257_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink200(
    .ins (cond_br257_falseOut),
    .ins_valid (cond_br257_falseOut_valid),
    .ins_ready (cond_br257_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(28)) cond_br258(
    .condition (fork78_outs_7),
    .condition_valid (fork78_outs_7_valid),
    .condition_ready (fork78_outs_7_ready),
    .data (constant544_outs),
    .data_valid (constant544_outs_valid),
    .data_ready (constant544_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br258_trueOut),
    .trueOut_valid (cond_br258_trueOut_valid),
    .trueOut_ready (cond_br258_trueOut_ready),
    .falseOut (cond_br258_falseOut),
    .falseOut_valid (cond_br258_falseOut_valid),
    .falseOut_ready (cond_br258_falseOut_ready)
  );

  sink #(.DATA_TYPE(28)) sink201(
    .ins (cond_br258_falseOut),
    .ins_valid (cond_br258_falseOut_valid),
    .ins_ready (cond_br258_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(28), .OUTPUT_TYPE(33)) extsi218(
    .ins (cond_br258_trueOut),
    .ins_valid (cond_br258_trueOut_valid),
    .ins_ready (cond_br258_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi218_outs),
    .outs_valid (extsi218_outs_valid),
    .outs_ready (extsi218_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br259(
    .condition (fork78_outs_3),
    .condition_valid (fork78_outs_3_valid),
    .condition_ready (fork78_outs_3_ready),
    .data (constant400_outs),
    .data_valid (constant400_outs_valid),
    .data_ready (constant400_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br259_trueOut),
    .trueOut_valid (cond_br259_trueOut_valid),
    .trueOut_ready (cond_br259_trueOut_ready),
    .falseOut (cond_br259_falseOut),
    .falseOut_valid (cond_br259_falseOut_valid),
    .falseOut_ready (cond_br259_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink202(
    .ins (cond_br259_falseOut),
    .ins_valid (cond_br259_falseOut_valid),
    .ins_ready (cond_br259_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(18)) cond_br260(
    .condition (fork78_outs_6),
    .condition_valid (fork78_outs_6_valid),
    .condition_ready (fork78_outs_6_ready),
    .data (constant545_outs),
    .data_valid (constant545_outs_valid),
    .data_ready (constant545_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br260_trueOut),
    .trueOut_valid (cond_br260_trueOut_valid),
    .trueOut_ready (cond_br260_trueOut_ready),
    .falseOut (cond_br260_falseOut),
    .falseOut_valid (cond_br260_falseOut_valid),
    .falseOut_ready (cond_br260_falseOut_ready)
  );

  sink #(.DATA_TYPE(18)) sink203(
    .ins (cond_br260_falseOut),
    .ins_valid (cond_br260_falseOut_valid),
    .ins_ready (cond_br260_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(18), .OUTPUT_TYPE(22)) extsi219(
    .ins (cond_br260_trueOut),
    .ins_valid (cond_br260_trueOut_valid),
    .ins_ready (cond_br260_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi219_outs),
    .outs_valid (extsi219_outs_valid),
    .outs_ready (extsi219_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br261(
    .condition (fork78_outs_2),
    .condition_valid (fork78_outs_2_valid),
    .condition_ready (fork78_outs_2_ready),
    .data (constant402_outs),
    .data_valid (constant402_outs_valid),
    .data_ready (constant402_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br261_trueOut),
    .trueOut_valid (cond_br261_trueOut_valid),
    .trueOut_ready (cond_br261_trueOut_ready),
    .falseOut (cond_br261_falseOut),
    .falseOut_valid (cond_br261_falseOut_valid),
    .falseOut_ready (cond_br261_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink204(
    .ins (cond_br261_falseOut),
    .ins_valid (cond_br261_falseOut_valid),
    .ins_ready (cond_br261_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br262(
    .condition (fork78_outs_5),
    .condition_valid (fork78_outs_5_valid),
    .condition_ready (fork78_outs_5_ready),
    .data (constant546_outs),
    .data_valid (constant546_outs_valid),
    .data_ready (constant546_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br262_trueOut),
    .trueOut_valid (cond_br262_trueOut_valid),
    .trueOut_ready (cond_br262_trueOut_ready),
    .falseOut (cond_br262_falseOut),
    .falseOut_valid (cond_br262_falseOut_valid),
    .falseOut_ready (cond_br262_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink205(
    .ins (cond_br262_falseOut),
    .ins_valid (cond_br262_falseOut_valid),
    .ins_ready (cond_br262_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(12)) extsi220(
    .ins (cond_br262_trueOut),
    .ins_valid (cond_br262_trueOut_valid),
    .ins_ready (cond_br262_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi220_outs),
    .outs_valid (extsi220_outs_valid),
    .outs_ready (extsi220_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer144(
    .ins (cond_br254_falseOut),
    .ins_valid (cond_br254_falseOut_valid),
    .ins_ready (cond_br254_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer144_outs),
    .outs_valid (buffer144_outs_valid),
    .outs_ready (buffer144_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer145(
    .ins (buffer144_outs),
    .ins_valid (buffer144_outs_valid),
    .ins_ready (buffer144_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer145_outs),
    .outs_valid (buffer145_outs_valid),
    .outs_ready (buffer145_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br263(
    .condition (fork78_outs_0),
    .condition_valid (fork78_outs_0_valid),
    .condition_ready (fork78_outs_0_ready),
    .data (buffer145_outs),
    .data_valid (buffer145_outs_valid),
    .data_ready (buffer145_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br263_trueOut),
    .trueOut_valid (cond_br263_trueOut_valid),
    .trueOut_ready (cond_br263_trueOut_ready),
    .falseOut (cond_br263_falseOut),
    .falseOut_valid (cond_br263_falseOut_valid),
    .falseOut_ready (cond_br263_falseOut_ready)
  );

  cond_br_dataless cond_br264(
    .condition (fork78_outs_1),
    .condition_valid (fork78_outs_1_valid),
    .condition_ready (fork78_outs_1_ready),
    .data_valid (fork77_outs_6_valid),
    .data_ready (fork77_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br264_trueOut_valid),
    .trueOut_ready (cond_br264_trueOut_ready),
    .falseOut_valid (cond_br264_falseOut_valid),
    .falseOut_ready (cond_br264_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br265(
    .condition (fork78_outs_8),
    .condition_valid (fork78_outs_8_valid),
    .condition_ready (fork78_outs_8_ready),
    .data (fork76_outs_1),
    .data_valid (fork76_outs_1_valid),
    .data_ready (fork76_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br265_trueOut),
    .trueOut_valid (cond_br265_trueOut_valid),
    .trueOut_ready (cond_br265_trueOut_ready),
    .falseOut (cond_br265_falseOut),
    .falseOut_valid (cond_br265_falseOut_valid),
    .falseOut_ready (cond_br265_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink206(
    .ins (cond_br265_trueOut),
    .ins_valid (cond_br265_trueOut_valid),
    .ins_ready (cond_br265_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer152(
    .ins (cond_br265_falseOut),
    .ins_valid (cond_br265_falseOut_valid),
    .ins_ready (cond_br265_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer152_outs),
    .outs_valid (buffer152_outs_valid),
    .outs_ready (buffer152_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer153(
    .ins (buffer152_outs),
    .ins_valid (buffer152_outs_valid),
    .ins_ready (buffer152_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer153_outs),
    .outs_valid (buffer153_outs_valid),
    .outs_ready (buffer153_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork79(
    .ins (buffer153_outs),
    .ins_valid (buffer153_outs_valid),
    .ins_ready (buffer153_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork79_outs_1, fork79_outs_0}),
    .outs_valid ({fork79_outs_1_valid, fork79_outs_0_valid}),
    .outs_ready ({fork79_outs_1_ready, fork79_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi221(
    .ins (fork79_outs_0),
    .ins_valid (fork79_outs_0_valid),
    .ins_ready (fork79_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi221_outs),
    .outs_valid (extsi221_outs_valid),
    .outs_ready (extsi221_outs_ready)
  );

  oehb_dataless buffer154(
    .ins_valid (cond_br264_falseOut_valid),
    .ins_ready (cond_br264_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer154_outs_valid),
    .outs_ready (buffer154_outs_ready)
  );

  tehb_dataless buffer155(
    .ins_valid (buffer154_outs_valid),
    .ins_ready (buffer154_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer155_outs_valid),
    .outs_ready (buffer155_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork80(
    .ins_valid (buffer155_outs_valid),
    .ins_ready (buffer155_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork80_outs_6_valid, fork80_outs_5_valid, fork80_outs_4_valid, fork80_outs_3_valid, fork80_outs_2_valid, fork80_outs_1_valid, fork80_outs_0_valid}),
    .outs_ready ({fork80_outs_6_ready, fork80_outs_5_ready, fork80_outs_4_ready, fork80_outs_3_ready, fork80_outs_2_ready, fork80_outs_1_ready, fork80_outs_0_ready})
  );

  handshake_constant_181 #(.DATA_WIDTH(37)) constant405(
    .ctrl_valid (fork80_outs_5_valid),
    .ctrl_ready (fork80_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant405_outs),
    .outs_valid (constant405_outs_valid),
    .outs_ready (constant405_outs_ready)
  );

  handshake_constant_182 #(.DATA_WIDTH(28)) constant548(
    .ctrl_valid (fork80_outs_2_valid),
    .ctrl_ready (fork80_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant548_outs),
    .outs_valid (constant548_outs_valid),
    .outs_ready (constant548_outs_ready)
  );

  handshake_constant_183 #(.DATA_WIDTH(27)) constant407(
    .ctrl_valid (fork80_outs_4_valid),
    .ctrl_ready (fork80_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant407_outs),
    .outs_valid (constant407_outs_valid),
    .outs_ready (constant407_outs_ready)
  );

  handshake_constant_184 #(.DATA_WIDTH(18)) constant549(
    .ctrl_valid (fork80_outs_1_valid),
    .ctrl_ready (fork80_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant549_outs),
    .outs_valid (constant549_outs_valid),
    .outs_ready (constant549_outs_ready)
  );

  handshake_constant_185 #(.DATA_WIDTH(17)) constant409(
    .ctrl_valid (fork80_outs_3_valid),
    .ctrl_ready (fork80_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant409_outs),
    .outs_valid (constant409_outs_valid),
    .outs_ready (constant409_outs_ready)
  );

  handshake_constant_186 #(.DATA_WIDTH(7)) constant550(
    .ctrl_valid (fork80_outs_0_valid),
    .ctrl_ready (fork80_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant550_outs),
    .outs_valid (constant550_outs_valid),
    .outs_ready (constant550_outs_ready)
  );

  source source27(
    .clk (clk),
    .rst (rst),
    .outs_valid (source27_outs_valid),
    .outs_ready (source27_outs_ready)
  );

  handshake_constant_187 #(.DATA_WIDTH(6)) constant551(
    .ctrl_valid (source27_outs_valid),
    .ctrl_ready (source27_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant551_outs),
    .outs_valid (constant551_outs_valid),
    .outs_ready (constant551_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi26(
    .lhs (extsi221_outs),
    .lhs_valid (extsi221_outs_valid),
    .lhs_ready (extsi221_outs_ready),
    .rhs (constant551_outs),
    .rhs_valid (constant551_outs_valid),
    .rhs_ready (constant551_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi26_result),
    .result_valid (cmpi26_result_valid),
    .result_ready (cmpi26_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork81(
    .ins (cmpi26_result),
    .ins_valid (cmpi26_result_valid),
    .ins_ready (cmpi26_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork81_outs_8, fork81_outs_7, fork81_outs_6, fork81_outs_5, fork81_outs_4, fork81_outs_3, fork81_outs_2, fork81_outs_1, fork81_outs_0}),
    .outs_valid ({fork81_outs_8_valid, fork81_outs_7_valid, fork81_outs_6_valid, fork81_outs_5_valid, fork81_outs_4_valid, fork81_outs_3_valid, fork81_outs_2_valid, fork81_outs_1_valid, fork81_outs_0_valid}),
    .outs_ready ({fork81_outs_8_ready, fork81_outs_7_ready, fork81_outs_6_ready, fork81_outs_5_ready, fork81_outs_4_ready, fork81_outs_3_ready, fork81_outs_2_ready, fork81_outs_1_ready, fork81_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br266(
    .condition (fork81_outs_4),
    .condition_valid (fork81_outs_4_valid),
    .condition_ready (fork81_outs_4_ready),
    .data (constant405_outs),
    .data_valid (constant405_outs_valid),
    .data_ready (constant405_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br266_trueOut),
    .trueOut_valid (cond_br266_trueOut_valid),
    .trueOut_ready (cond_br266_trueOut_ready),
    .falseOut (cond_br266_falseOut),
    .falseOut_valid (cond_br266_falseOut_valid),
    .falseOut_ready (cond_br266_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink208(
    .ins (cond_br266_falseOut),
    .ins_valid (cond_br266_falseOut_valid),
    .ins_ready (cond_br266_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(28)) cond_br267(
    .condition (fork81_outs_7),
    .condition_valid (fork81_outs_7_valid),
    .condition_ready (fork81_outs_7_ready),
    .data (constant548_outs),
    .data_valid (constant548_outs_valid),
    .data_ready (constant548_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br267_trueOut),
    .trueOut_valid (cond_br267_trueOut_valid),
    .trueOut_ready (cond_br267_trueOut_ready),
    .falseOut (cond_br267_falseOut),
    .falseOut_valid (cond_br267_falseOut_valid),
    .falseOut_ready (cond_br267_falseOut_ready)
  );

  sink #(.DATA_TYPE(28)) sink209(
    .ins (cond_br267_falseOut),
    .ins_valid (cond_br267_falseOut_valid),
    .ins_ready (cond_br267_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(28), .OUTPUT_TYPE(33)) extsi222(
    .ins (cond_br267_trueOut),
    .ins_valid (cond_br267_trueOut_valid),
    .ins_ready (cond_br267_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi222_outs),
    .outs_valid (extsi222_outs_valid),
    .outs_ready (extsi222_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br268(
    .condition (fork81_outs_3),
    .condition_valid (fork81_outs_3_valid),
    .condition_ready (fork81_outs_3_ready),
    .data (constant407_outs),
    .data_valid (constant407_outs_valid),
    .data_ready (constant407_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br268_trueOut),
    .trueOut_valid (cond_br268_trueOut_valid),
    .trueOut_ready (cond_br268_trueOut_ready),
    .falseOut (cond_br268_falseOut),
    .falseOut_valid (cond_br268_falseOut_valid),
    .falseOut_ready (cond_br268_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink210(
    .ins (cond_br268_falseOut),
    .ins_valid (cond_br268_falseOut_valid),
    .ins_ready (cond_br268_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(18)) cond_br269(
    .condition (fork81_outs_6),
    .condition_valid (fork81_outs_6_valid),
    .condition_ready (fork81_outs_6_ready),
    .data (constant549_outs),
    .data_valid (constant549_outs_valid),
    .data_ready (constant549_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br269_trueOut),
    .trueOut_valid (cond_br269_trueOut_valid),
    .trueOut_ready (cond_br269_trueOut_ready),
    .falseOut (cond_br269_falseOut),
    .falseOut_valid (cond_br269_falseOut_valid),
    .falseOut_ready (cond_br269_falseOut_ready)
  );

  sink #(.DATA_TYPE(18)) sink211(
    .ins (cond_br269_falseOut),
    .ins_valid (cond_br269_falseOut_valid),
    .ins_ready (cond_br269_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(18), .OUTPUT_TYPE(22)) extsi223(
    .ins (cond_br269_trueOut),
    .ins_valid (cond_br269_trueOut_valid),
    .ins_ready (cond_br269_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi223_outs),
    .outs_valid (extsi223_outs_valid),
    .outs_ready (extsi223_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br270(
    .condition (fork81_outs_2),
    .condition_valid (fork81_outs_2_valid),
    .condition_ready (fork81_outs_2_ready),
    .data (constant409_outs),
    .data_valid (constant409_outs_valid),
    .data_ready (constant409_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br270_trueOut),
    .trueOut_valid (cond_br270_trueOut_valid),
    .trueOut_ready (cond_br270_trueOut_ready),
    .falseOut (cond_br270_falseOut),
    .falseOut_valid (cond_br270_falseOut_valid),
    .falseOut_ready (cond_br270_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink212(
    .ins (cond_br270_falseOut),
    .ins_valid (cond_br270_falseOut_valid),
    .ins_ready (cond_br270_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br271(
    .condition (fork81_outs_5),
    .condition_valid (fork81_outs_5_valid),
    .condition_ready (fork81_outs_5_ready),
    .data (constant550_outs),
    .data_valid (constant550_outs_valid),
    .data_ready (constant550_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br271_trueOut),
    .trueOut_valid (cond_br271_trueOut_valid),
    .trueOut_ready (cond_br271_trueOut_ready),
    .falseOut (cond_br271_falseOut),
    .falseOut_valid (cond_br271_falseOut_valid),
    .falseOut_ready (cond_br271_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink213(
    .ins (cond_br271_falseOut),
    .ins_valid (cond_br271_falseOut_valid),
    .ins_ready (cond_br271_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(12)) extsi224(
    .ins (cond_br271_trueOut),
    .ins_valid (cond_br271_trueOut_valid),
    .ins_ready (cond_br271_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi224_outs),
    .outs_valid (extsi224_outs_valid),
    .outs_ready (extsi224_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer150(
    .ins (cond_br263_falseOut),
    .ins_valid (cond_br263_falseOut_valid),
    .ins_ready (cond_br263_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer150_outs),
    .outs_valid (buffer150_outs_valid),
    .outs_ready (buffer150_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer151(
    .ins (buffer150_outs),
    .ins_valid (buffer150_outs_valid),
    .ins_ready (buffer150_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer151_outs),
    .outs_valid (buffer151_outs_valid),
    .outs_ready (buffer151_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br272(
    .condition (fork81_outs_0),
    .condition_valid (fork81_outs_0_valid),
    .condition_ready (fork81_outs_0_ready),
    .data (buffer151_outs),
    .data_valid (buffer151_outs_valid),
    .data_ready (buffer151_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br272_trueOut),
    .trueOut_valid (cond_br272_trueOut_valid),
    .trueOut_ready (cond_br272_trueOut_ready),
    .falseOut (cond_br272_falseOut),
    .falseOut_valid (cond_br272_falseOut_valid),
    .falseOut_ready (cond_br272_falseOut_ready)
  );

  cond_br_dataless cond_br273(
    .condition (fork81_outs_1),
    .condition_valid (fork81_outs_1_valid),
    .condition_ready (fork81_outs_1_ready),
    .data_valid (fork80_outs_6_valid),
    .data_ready (fork80_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br273_trueOut_valid),
    .trueOut_ready (cond_br273_trueOut_ready),
    .falseOut_valid (cond_br273_falseOut_valid),
    .falseOut_ready (cond_br273_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br274(
    .condition (fork81_outs_8),
    .condition_valid (fork81_outs_8_valid),
    .condition_ready (fork81_outs_8_ready),
    .data (fork79_outs_1),
    .data_valid (fork79_outs_1_valid),
    .data_ready (fork79_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br274_trueOut),
    .trueOut_valid (cond_br274_trueOut_valid),
    .trueOut_ready (cond_br274_trueOut_ready),
    .falseOut (cond_br274_falseOut),
    .falseOut_valid (cond_br274_falseOut_valid),
    .falseOut_ready (cond_br274_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink214(
    .ins (cond_br274_trueOut),
    .ins_valid (cond_br274_trueOut_valid),
    .ins_ready (cond_br274_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer158(
    .ins (cond_br274_falseOut),
    .ins_valid (cond_br274_falseOut_valid),
    .ins_ready (cond_br274_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer158_outs),
    .outs_valid (buffer158_outs_valid),
    .outs_ready (buffer158_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer159(
    .ins (buffer158_outs),
    .ins_valid (buffer158_outs_valid),
    .ins_ready (buffer158_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer159_outs),
    .outs_valid (buffer159_outs_valid),
    .outs_ready (buffer159_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork82(
    .ins (buffer159_outs),
    .ins_valid (buffer159_outs_valid),
    .ins_ready (buffer159_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork82_outs_1, fork82_outs_0}),
    .outs_valid ({fork82_outs_1_valid, fork82_outs_0_valid}),
    .outs_ready ({fork82_outs_1_ready, fork82_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi225(
    .ins (fork82_outs_0),
    .ins_valid (fork82_outs_0_valid),
    .ins_ready (fork82_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi225_outs),
    .outs_valid (extsi225_outs_valid),
    .outs_ready (extsi225_outs_ready)
  );

  oehb_dataless buffer160(
    .ins_valid (cond_br273_falseOut_valid),
    .ins_ready (cond_br273_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer160_outs_valid),
    .outs_ready (buffer160_outs_ready)
  );

  tehb_dataless buffer161(
    .ins_valid (buffer160_outs_valid),
    .ins_ready (buffer160_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer161_outs_valid),
    .outs_ready (buffer161_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork83(
    .ins_valid (buffer161_outs_valid),
    .ins_ready (buffer161_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork83_outs_6_valid, fork83_outs_5_valid, fork83_outs_4_valid, fork83_outs_3_valid, fork83_outs_2_valid, fork83_outs_1_valid, fork83_outs_0_valid}),
    .outs_ready ({fork83_outs_6_ready, fork83_outs_5_ready, fork83_outs_4_ready, fork83_outs_3_ready, fork83_outs_2_ready, fork83_outs_1_ready, fork83_outs_0_ready})
  );

  handshake_constant_188 #(.DATA_WIDTH(37)) constant412(
    .ctrl_valid (fork83_outs_5_valid),
    .ctrl_ready (fork83_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant412_outs),
    .outs_valid (constant412_outs_valid),
    .outs_ready (constant412_outs_ready)
  );

  handshake_constant_189 #(.DATA_WIDTH(27)) constant552(
    .ctrl_valid (fork83_outs_2_valid),
    .ctrl_ready (fork83_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant552_outs),
    .outs_valid (constant552_outs_valid),
    .outs_ready (constant552_outs_ready)
  );

  handshake_constant_190 #(.DATA_WIDTH(27)) constant414(
    .ctrl_valid (fork83_outs_4_valid),
    .ctrl_ready (fork83_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant414_outs),
    .outs_valid (constant414_outs_valid),
    .outs_ready (constant414_outs_ready)
  );

  handshake_constant_191 #(.DATA_WIDTH(18)) constant553(
    .ctrl_valid (fork83_outs_1_valid),
    .ctrl_ready (fork83_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant553_outs),
    .outs_valid (constant553_outs_valid),
    .outs_ready (constant553_outs_ready)
  );

  handshake_constant_192 #(.DATA_WIDTH(17)) constant416(
    .ctrl_valid (fork83_outs_3_valid),
    .ctrl_ready (fork83_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant416_outs),
    .outs_valid (constant416_outs_valid),
    .outs_ready (constant416_outs_ready)
  );

  handshake_constant_193 #(.DATA_WIDTH(7)) constant554(
    .ctrl_valid (fork83_outs_0_valid),
    .ctrl_ready (fork83_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant554_outs),
    .outs_valid (constant554_outs_valid),
    .outs_ready (constant554_outs_ready)
  );

  source source28(
    .clk (clk),
    .rst (rst),
    .outs_valid (source28_outs_valid),
    .outs_ready (source28_outs_ready)
  );

  handshake_constant_124 #(.DATA_WIDTH(6)) constant555(
    .ctrl_valid (source28_outs_valid),
    .ctrl_ready (source28_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant555_outs),
    .outs_valid (constant555_outs_valid),
    .outs_ready (constant555_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi27(
    .lhs (extsi225_outs),
    .lhs_valid (extsi225_outs_valid),
    .lhs_ready (extsi225_outs_ready),
    .rhs (constant555_outs),
    .rhs_valid (constant555_outs_valid),
    .rhs_ready (constant555_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi27_result),
    .result_valid (cmpi27_result_valid),
    .result_ready (cmpi27_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork84(
    .ins (cmpi27_result),
    .ins_valid (cmpi27_result_valid),
    .ins_ready (cmpi27_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork84_outs_8, fork84_outs_7, fork84_outs_6, fork84_outs_5, fork84_outs_4, fork84_outs_3, fork84_outs_2, fork84_outs_1, fork84_outs_0}),
    .outs_valid ({fork84_outs_8_valid, fork84_outs_7_valid, fork84_outs_6_valid, fork84_outs_5_valid, fork84_outs_4_valid, fork84_outs_3_valid, fork84_outs_2_valid, fork84_outs_1_valid, fork84_outs_0_valid}),
    .outs_ready ({fork84_outs_8_ready, fork84_outs_7_ready, fork84_outs_6_ready, fork84_outs_5_ready, fork84_outs_4_ready, fork84_outs_3_ready, fork84_outs_2_ready, fork84_outs_1_ready, fork84_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br275(
    .condition (fork84_outs_4),
    .condition_valid (fork84_outs_4_valid),
    .condition_ready (fork84_outs_4_ready),
    .data (constant412_outs),
    .data_valid (constant412_outs_valid),
    .data_ready (constant412_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br275_trueOut),
    .trueOut_valid (cond_br275_trueOut_valid),
    .trueOut_ready (cond_br275_trueOut_ready),
    .falseOut (cond_br275_falseOut),
    .falseOut_valid (cond_br275_falseOut_valid),
    .falseOut_ready (cond_br275_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink216(
    .ins (cond_br275_falseOut),
    .ins_valid (cond_br275_falseOut_valid),
    .ins_ready (cond_br275_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br276(
    .condition (fork84_outs_7),
    .condition_valid (fork84_outs_7_valid),
    .condition_ready (fork84_outs_7_ready),
    .data (constant552_outs),
    .data_valid (constant552_outs_valid),
    .data_ready (constant552_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br276_trueOut),
    .trueOut_valid (cond_br276_trueOut_valid),
    .trueOut_ready (cond_br276_trueOut_ready),
    .falseOut (cond_br276_falseOut),
    .falseOut_valid (cond_br276_falseOut_valid),
    .falseOut_ready (cond_br276_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink217(
    .ins (cond_br276_falseOut),
    .ins_valid (cond_br276_falseOut_valid),
    .ins_ready (cond_br276_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(27), .OUTPUT_TYPE(33)) extsi226(
    .ins (cond_br276_trueOut),
    .ins_valid (cond_br276_trueOut_valid),
    .ins_ready (cond_br276_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi226_outs),
    .outs_valid (extsi226_outs_valid),
    .outs_ready (extsi226_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br277(
    .condition (fork84_outs_3),
    .condition_valid (fork84_outs_3_valid),
    .condition_ready (fork84_outs_3_ready),
    .data (constant414_outs),
    .data_valid (constant414_outs_valid),
    .data_ready (constant414_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br277_trueOut),
    .trueOut_valid (cond_br277_trueOut_valid),
    .trueOut_ready (cond_br277_trueOut_ready),
    .falseOut (cond_br277_falseOut),
    .falseOut_valid (cond_br277_falseOut_valid),
    .falseOut_ready (cond_br277_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink218(
    .ins (cond_br277_falseOut),
    .ins_valid (cond_br277_falseOut_valid),
    .ins_ready (cond_br277_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(18)) cond_br278(
    .condition (fork84_outs_6),
    .condition_valid (fork84_outs_6_valid),
    .condition_ready (fork84_outs_6_ready),
    .data (constant553_outs),
    .data_valid (constant553_outs_valid),
    .data_ready (constant553_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br278_trueOut),
    .trueOut_valid (cond_br278_trueOut_valid),
    .trueOut_ready (cond_br278_trueOut_ready),
    .falseOut (cond_br278_falseOut),
    .falseOut_valid (cond_br278_falseOut_valid),
    .falseOut_ready (cond_br278_falseOut_ready)
  );

  sink #(.DATA_TYPE(18)) sink219(
    .ins (cond_br278_falseOut),
    .ins_valid (cond_br278_falseOut_valid),
    .ins_ready (cond_br278_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(18), .OUTPUT_TYPE(22)) extsi227(
    .ins (cond_br278_trueOut),
    .ins_valid (cond_br278_trueOut_valid),
    .ins_ready (cond_br278_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi227_outs),
    .outs_valid (extsi227_outs_valid),
    .outs_ready (extsi227_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br279(
    .condition (fork84_outs_2),
    .condition_valid (fork84_outs_2_valid),
    .condition_ready (fork84_outs_2_ready),
    .data (constant416_outs),
    .data_valid (constant416_outs_valid),
    .data_ready (constant416_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br279_trueOut),
    .trueOut_valid (cond_br279_trueOut_valid),
    .trueOut_ready (cond_br279_trueOut_ready),
    .falseOut (cond_br279_falseOut),
    .falseOut_valid (cond_br279_falseOut_valid),
    .falseOut_ready (cond_br279_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink220(
    .ins (cond_br279_falseOut),
    .ins_valid (cond_br279_falseOut_valid),
    .ins_ready (cond_br279_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(7)) cond_br280(
    .condition (fork84_outs_5),
    .condition_valid (fork84_outs_5_valid),
    .condition_ready (fork84_outs_5_ready),
    .data (constant554_outs),
    .data_valid (constant554_outs_valid),
    .data_ready (constant554_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br280_trueOut),
    .trueOut_valid (cond_br280_trueOut_valid),
    .trueOut_ready (cond_br280_trueOut_ready),
    .falseOut (cond_br280_falseOut),
    .falseOut_valid (cond_br280_falseOut_valid),
    .falseOut_ready (cond_br280_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink221(
    .ins (cond_br280_falseOut),
    .ins_valid (cond_br280_falseOut_valid),
    .ins_ready (cond_br280_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(12)) extsi228(
    .ins (cond_br280_trueOut),
    .ins_valid (cond_br280_trueOut_valid),
    .ins_ready (cond_br280_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi228_outs),
    .outs_valid (extsi228_outs_valid),
    .outs_ready (extsi228_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer156(
    .ins (cond_br272_falseOut),
    .ins_valid (cond_br272_falseOut_valid),
    .ins_ready (cond_br272_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer156_outs),
    .outs_valid (buffer156_outs_valid),
    .outs_ready (buffer156_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer157(
    .ins (buffer156_outs),
    .ins_valid (buffer156_outs_valid),
    .ins_ready (buffer156_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer157_outs),
    .outs_valid (buffer157_outs_valid),
    .outs_ready (buffer157_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br281(
    .condition (fork84_outs_0),
    .condition_valid (fork84_outs_0_valid),
    .condition_ready (fork84_outs_0_ready),
    .data (buffer157_outs),
    .data_valid (buffer157_outs_valid),
    .data_ready (buffer157_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br281_trueOut),
    .trueOut_valid (cond_br281_trueOut_valid),
    .trueOut_ready (cond_br281_trueOut_ready),
    .falseOut (cond_br281_falseOut),
    .falseOut_valid (cond_br281_falseOut_valid),
    .falseOut_ready (cond_br281_falseOut_ready)
  );

  cond_br_dataless cond_br282(
    .condition (fork84_outs_1),
    .condition_valid (fork84_outs_1_valid),
    .condition_ready (fork84_outs_1_ready),
    .data_valid (fork83_outs_6_valid),
    .data_ready (fork83_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br282_trueOut_valid),
    .trueOut_ready (cond_br282_trueOut_ready),
    .falseOut_valid (cond_br282_falseOut_valid),
    .falseOut_ready (cond_br282_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br283(
    .condition (fork84_outs_8),
    .condition_valid (fork84_outs_8_valid),
    .condition_ready (fork84_outs_8_ready),
    .data (fork82_outs_1),
    .data_valid (fork82_outs_1_valid),
    .data_ready (fork82_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br283_trueOut),
    .trueOut_valid (cond_br283_trueOut_valid),
    .trueOut_ready (cond_br283_trueOut_ready),
    .falseOut (cond_br283_falseOut),
    .falseOut_valid (cond_br283_falseOut_valid),
    .falseOut_ready (cond_br283_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink222(
    .ins (cond_br283_trueOut),
    .ins_valid (cond_br283_trueOut_valid),
    .ins_ready (cond_br283_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer164(
    .ins (cond_br283_falseOut),
    .ins_valid (cond_br283_falseOut_valid),
    .ins_ready (cond_br283_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer164_outs),
    .outs_valid (buffer164_outs_valid),
    .outs_ready (buffer164_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer165(
    .ins (buffer164_outs),
    .ins_valid (buffer164_outs_valid),
    .ins_ready (buffer164_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer165_outs),
    .outs_valid (buffer165_outs_valid),
    .outs_ready (buffer165_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork85(
    .ins (buffer165_outs),
    .ins_valid (buffer165_outs_valid),
    .ins_ready (buffer165_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork85_outs_1, fork85_outs_0}),
    .outs_valid ({fork85_outs_1_valid, fork85_outs_0_valid}),
    .outs_ready ({fork85_outs_1_ready, fork85_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi229(
    .ins (fork85_outs_0),
    .ins_valid (fork85_outs_0_valid),
    .ins_ready (fork85_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi229_outs),
    .outs_valid (extsi229_outs_valid),
    .outs_ready (extsi229_outs_ready)
  );

  oehb_dataless buffer166(
    .ins_valid (cond_br282_falseOut_valid),
    .ins_ready (cond_br282_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer166_outs_valid),
    .outs_ready (buffer166_outs_ready)
  );

  tehb_dataless buffer167(
    .ins_valid (buffer166_outs_valid),
    .ins_ready (buffer166_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer167_outs_valid),
    .outs_ready (buffer167_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork86(
    .ins_valid (buffer167_outs_valid),
    .ins_ready (buffer167_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork86_outs_6_valid, fork86_outs_5_valid, fork86_outs_4_valid, fork86_outs_3_valid, fork86_outs_2_valid, fork86_outs_1_valid, fork86_outs_0_valid}),
    .outs_ready ({fork86_outs_6_ready, fork86_outs_5_ready, fork86_outs_4_ready, fork86_outs_3_ready, fork86_outs_2_ready, fork86_outs_1_ready, fork86_outs_0_ready})
  );

  handshake_constant_194 #(.DATA_WIDTH(37)) constant419(
    .ctrl_valid (fork86_outs_5_valid),
    .ctrl_ready (fork86_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant419_outs),
    .outs_valid (constant419_outs_valid),
    .outs_ready (constant419_outs_ready)
  );

  handshake_constant_195 #(.DATA_WIDTH(27)) constant556(
    .ctrl_valid (fork86_outs_2_valid),
    .ctrl_ready (fork86_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant556_outs),
    .outs_valid (constant556_outs_valid),
    .outs_ready (constant556_outs_ready)
  );

  handshake_constant_196 #(.DATA_WIDTH(27)) constant421(
    .ctrl_valid (fork86_outs_4_valid),
    .ctrl_ready (fork86_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant421_outs),
    .outs_valid (constant421_outs_valid),
    .outs_ready (constant421_outs_ready)
  );

  handshake_constant_197 #(.DATA_WIDTH(18)) constant557(
    .ctrl_valid (fork86_outs_1_valid),
    .ctrl_ready (fork86_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant557_outs),
    .outs_valid (constant557_outs_valid),
    .outs_ready (constant557_outs_ready)
  );

  handshake_constant_198 #(.DATA_WIDTH(17)) constant423(
    .ctrl_valid (fork86_outs_3_valid),
    .ctrl_ready (fork86_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant423_outs),
    .outs_valid (constant423_outs_valid),
    .outs_ready (constant423_outs_ready)
  );

  handshake_constant_199 #(.DATA_WIDTH(6)) constant558(
    .ctrl_valid (fork86_outs_0_valid),
    .ctrl_ready (fork86_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant558_outs),
    .outs_valid (constant558_outs_valid),
    .outs_ready (constant558_outs_ready)
  );

  source source29(
    .clk (clk),
    .rst (rst),
    .outs_valid (source29_outs_valid),
    .outs_ready (source29_outs_ready)
  );

  handshake_constant_200 #(.DATA_WIDTH(6)) constant559(
    .ctrl_valid (source29_outs_valid),
    .ctrl_ready (source29_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant559_outs),
    .outs_valid (constant559_outs_valid),
    .outs_ready (constant559_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi28(
    .lhs (extsi229_outs),
    .lhs_valid (extsi229_outs_valid),
    .lhs_ready (extsi229_outs_ready),
    .rhs (constant559_outs),
    .rhs_valid (constant559_outs_valid),
    .rhs_ready (constant559_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi28_result),
    .result_valid (cmpi28_result_valid),
    .result_ready (cmpi28_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork87(
    .ins (cmpi28_result),
    .ins_valid (cmpi28_result_valid),
    .ins_ready (cmpi28_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork87_outs_8, fork87_outs_7, fork87_outs_6, fork87_outs_5, fork87_outs_4, fork87_outs_3, fork87_outs_2, fork87_outs_1, fork87_outs_0}),
    .outs_valid ({fork87_outs_8_valid, fork87_outs_7_valid, fork87_outs_6_valid, fork87_outs_5_valid, fork87_outs_4_valid, fork87_outs_3_valid, fork87_outs_2_valid, fork87_outs_1_valid, fork87_outs_0_valid}),
    .outs_ready ({fork87_outs_8_ready, fork87_outs_7_ready, fork87_outs_6_ready, fork87_outs_5_ready, fork87_outs_4_ready, fork87_outs_3_ready, fork87_outs_2_ready, fork87_outs_1_ready, fork87_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br284(
    .condition (fork87_outs_4),
    .condition_valid (fork87_outs_4_valid),
    .condition_ready (fork87_outs_4_ready),
    .data (constant419_outs),
    .data_valid (constant419_outs_valid),
    .data_ready (constant419_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br284_trueOut),
    .trueOut_valid (cond_br284_trueOut_valid),
    .trueOut_ready (cond_br284_trueOut_ready),
    .falseOut (cond_br284_falseOut),
    .falseOut_valid (cond_br284_falseOut_valid),
    .falseOut_ready (cond_br284_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink224(
    .ins (cond_br284_falseOut),
    .ins_valid (cond_br284_falseOut_valid),
    .ins_ready (cond_br284_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br285(
    .condition (fork87_outs_7),
    .condition_valid (fork87_outs_7_valid),
    .condition_ready (fork87_outs_7_ready),
    .data (constant556_outs),
    .data_valid (constant556_outs_valid),
    .data_ready (constant556_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br285_trueOut),
    .trueOut_valid (cond_br285_trueOut_valid),
    .trueOut_ready (cond_br285_trueOut_ready),
    .falseOut (cond_br285_falseOut),
    .falseOut_valid (cond_br285_falseOut_valid),
    .falseOut_ready (cond_br285_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink225(
    .ins (cond_br285_falseOut),
    .ins_valid (cond_br285_falseOut_valid),
    .ins_ready (cond_br285_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(27), .OUTPUT_TYPE(33)) extsi230(
    .ins (cond_br285_trueOut),
    .ins_valid (cond_br285_trueOut_valid),
    .ins_ready (cond_br285_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi230_outs),
    .outs_valid (extsi230_outs_valid),
    .outs_ready (extsi230_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br286(
    .condition (fork87_outs_3),
    .condition_valid (fork87_outs_3_valid),
    .condition_ready (fork87_outs_3_ready),
    .data (constant421_outs),
    .data_valid (constant421_outs_valid),
    .data_ready (constant421_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br286_trueOut),
    .trueOut_valid (cond_br286_trueOut_valid),
    .trueOut_ready (cond_br286_trueOut_ready),
    .falseOut (cond_br286_falseOut),
    .falseOut_valid (cond_br286_falseOut_valid),
    .falseOut_ready (cond_br286_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink226(
    .ins (cond_br286_falseOut),
    .ins_valid (cond_br286_falseOut_valid),
    .ins_ready (cond_br286_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(18)) cond_br287(
    .condition (fork87_outs_6),
    .condition_valid (fork87_outs_6_valid),
    .condition_ready (fork87_outs_6_ready),
    .data (constant557_outs),
    .data_valid (constant557_outs_valid),
    .data_ready (constant557_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br287_trueOut),
    .trueOut_valid (cond_br287_trueOut_valid),
    .trueOut_ready (cond_br287_trueOut_ready),
    .falseOut (cond_br287_falseOut),
    .falseOut_valid (cond_br287_falseOut_valid),
    .falseOut_ready (cond_br287_falseOut_ready)
  );

  sink #(.DATA_TYPE(18)) sink227(
    .ins (cond_br287_falseOut),
    .ins_valid (cond_br287_falseOut_valid),
    .ins_ready (cond_br287_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(18), .OUTPUT_TYPE(22)) extsi231(
    .ins (cond_br287_trueOut),
    .ins_valid (cond_br287_trueOut_valid),
    .ins_ready (cond_br287_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi231_outs),
    .outs_valid (extsi231_outs_valid),
    .outs_ready (extsi231_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br288(
    .condition (fork87_outs_2),
    .condition_valid (fork87_outs_2_valid),
    .condition_ready (fork87_outs_2_ready),
    .data (constant423_outs),
    .data_valid (constant423_outs_valid),
    .data_ready (constant423_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br288_trueOut),
    .trueOut_valid (cond_br288_trueOut_valid),
    .trueOut_ready (cond_br288_trueOut_ready),
    .falseOut (cond_br288_falseOut),
    .falseOut_valid (cond_br288_falseOut_valid),
    .falseOut_ready (cond_br288_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink228(
    .ins (cond_br288_falseOut),
    .ins_valid (cond_br288_falseOut_valid),
    .ins_ready (cond_br288_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(6)) cond_br289(
    .condition (fork87_outs_5),
    .condition_valid (fork87_outs_5_valid),
    .condition_ready (fork87_outs_5_ready),
    .data (constant558_outs),
    .data_valid (constant558_outs_valid),
    .data_ready (constant558_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br289_trueOut),
    .trueOut_valid (cond_br289_trueOut_valid),
    .trueOut_ready (cond_br289_trueOut_ready),
    .falseOut (cond_br289_falseOut),
    .falseOut_valid (cond_br289_falseOut_valid),
    .falseOut_ready (cond_br289_falseOut_ready)
  );

  sink #(.DATA_TYPE(6)) sink229(
    .ins (cond_br289_falseOut),
    .ins_valid (cond_br289_falseOut_valid),
    .ins_ready (cond_br289_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(12)) extsi232(
    .ins (cond_br289_trueOut),
    .ins_valid (cond_br289_trueOut_valid),
    .ins_ready (cond_br289_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi232_outs),
    .outs_valid (extsi232_outs_valid),
    .outs_ready (extsi232_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer162(
    .ins (cond_br281_falseOut),
    .ins_valid (cond_br281_falseOut_valid),
    .ins_ready (cond_br281_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer162_outs),
    .outs_valid (buffer162_outs_valid),
    .outs_ready (buffer162_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer163(
    .ins (buffer162_outs),
    .ins_valid (buffer162_outs_valid),
    .ins_ready (buffer162_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer163_outs),
    .outs_valid (buffer163_outs_valid),
    .outs_ready (buffer163_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br290(
    .condition (fork87_outs_0),
    .condition_valid (fork87_outs_0_valid),
    .condition_ready (fork87_outs_0_ready),
    .data (buffer163_outs),
    .data_valid (buffer163_outs_valid),
    .data_ready (buffer163_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br290_trueOut),
    .trueOut_valid (cond_br290_trueOut_valid),
    .trueOut_ready (cond_br290_trueOut_ready),
    .falseOut (cond_br290_falseOut),
    .falseOut_valid (cond_br290_falseOut_valid),
    .falseOut_ready (cond_br290_falseOut_ready)
  );

  cond_br_dataless cond_br291(
    .condition (fork87_outs_1),
    .condition_valid (fork87_outs_1_valid),
    .condition_ready (fork87_outs_1_ready),
    .data_valid (fork86_outs_6_valid),
    .data_ready (fork86_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br291_trueOut_valid),
    .trueOut_ready (cond_br291_trueOut_ready),
    .falseOut_valid (cond_br291_falseOut_valid),
    .falseOut_ready (cond_br291_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br292(
    .condition (fork87_outs_8),
    .condition_valid (fork87_outs_8_valid),
    .condition_ready (fork87_outs_8_ready),
    .data (fork85_outs_1),
    .data_valid (fork85_outs_1_valid),
    .data_ready (fork85_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br292_trueOut),
    .trueOut_valid (cond_br292_trueOut_valid),
    .trueOut_ready (cond_br292_trueOut_ready),
    .falseOut (cond_br292_falseOut),
    .falseOut_valid (cond_br292_falseOut_valid),
    .falseOut_ready (cond_br292_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink230(
    .ins (cond_br292_trueOut),
    .ins_valid (cond_br292_trueOut_valid),
    .ins_ready (cond_br292_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer170(
    .ins (cond_br292_falseOut),
    .ins_valid (cond_br292_falseOut_valid),
    .ins_ready (cond_br292_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer170_outs),
    .outs_valid (buffer170_outs_valid),
    .outs_ready (buffer170_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer171(
    .ins (buffer170_outs),
    .ins_valid (buffer170_outs_valid),
    .ins_ready (buffer170_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer171_outs),
    .outs_valid (buffer171_outs_valid),
    .outs_ready (buffer171_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork88(
    .ins (buffer171_outs),
    .ins_valid (buffer171_outs_valid),
    .ins_ready (buffer171_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork88_outs_1, fork88_outs_0}),
    .outs_valid ({fork88_outs_1_valid, fork88_outs_0_valid}),
    .outs_ready ({fork88_outs_1_ready, fork88_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi233(
    .ins (fork88_outs_0),
    .ins_valid (fork88_outs_0_valid),
    .ins_ready (fork88_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi233_outs),
    .outs_valid (extsi233_outs_valid),
    .outs_ready (extsi233_outs_ready)
  );

  oehb_dataless buffer172(
    .ins_valid (cond_br291_falseOut_valid),
    .ins_ready (cond_br291_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer172_outs_valid),
    .outs_ready (buffer172_outs_ready)
  );

  tehb_dataless buffer173(
    .ins_valid (buffer172_outs_valid),
    .ins_ready (buffer172_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer173_outs_valid),
    .outs_ready (buffer173_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork89(
    .ins_valid (buffer173_outs_valid),
    .ins_ready (buffer173_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork89_outs_6_valid, fork89_outs_5_valid, fork89_outs_4_valid, fork89_outs_3_valid, fork89_outs_2_valid, fork89_outs_1_valid, fork89_outs_0_valid}),
    .outs_ready ({fork89_outs_6_ready, fork89_outs_5_ready, fork89_outs_4_ready, fork89_outs_3_ready, fork89_outs_2_ready, fork89_outs_1_ready, fork89_outs_0_ready})
  );

  handshake_constant_201 #(.DATA_WIDTH(37)) constant426(
    .ctrl_valid (fork89_outs_5_valid),
    .ctrl_ready (fork89_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant426_outs),
    .outs_valid (constant426_outs_valid),
    .outs_ready (constant426_outs_ready)
  );

  handshake_constant_202 #(.DATA_WIDTH(27)) constant560(
    .ctrl_valid (fork89_outs_2_valid),
    .ctrl_ready (fork89_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant560_outs),
    .outs_valid (constant560_outs_valid),
    .outs_ready (constant560_outs_ready)
  );

  handshake_constant_203 #(.DATA_WIDTH(27)) constant428(
    .ctrl_valid (fork89_outs_4_valid),
    .ctrl_ready (fork89_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant428_outs),
    .outs_valid (constant428_outs_valid),
    .outs_ready (constant428_outs_ready)
  );

  handshake_constant_204 #(.DATA_WIDTH(17)) constant561(
    .ctrl_valid (fork89_outs_1_valid),
    .ctrl_ready (fork89_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant561_outs),
    .outs_valid (constant561_outs_valid),
    .outs_ready (constant561_outs_ready)
  );

  handshake_constant_205 #(.DATA_WIDTH(17)) constant430(
    .ctrl_valid (fork89_outs_3_valid),
    .ctrl_ready (fork89_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant430_outs),
    .outs_valid (constant430_outs_valid),
    .outs_ready (constant430_outs_ready)
  );

  handshake_constant_166 #(.DATA_WIDTH(6)) constant562(
    .ctrl_valid (fork89_outs_0_valid),
    .ctrl_ready (fork89_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant562_outs),
    .outs_valid (constant562_outs_valid),
    .outs_ready (constant562_outs_ready)
  );

  source source30(
    .clk (clk),
    .rst (rst),
    .outs_valid (source30_outs_valid),
    .outs_ready (source30_outs_ready)
  );

  handshake_constant_206 #(.DATA_WIDTH(6)) constant563(
    .ctrl_valid (source30_outs_valid),
    .ctrl_ready (source30_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant563_outs),
    .outs_valid (constant563_outs_valid),
    .outs_ready (constant563_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi29(
    .lhs (extsi233_outs),
    .lhs_valid (extsi233_outs_valid),
    .lhs_ready (extsi233_outs_ready),
    .rhs (constant563_outs),
    .rhs_valid (constant563_outs_valid),
    .rhs_ready (constant563_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi29_result),
    .result_valid (cmpi29_result_valid),
    .result_ready (cmpi29_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork90(
    .ins (cmpi29_result),
    .ins_valid (cmpi29_result_valid),
    .ins_ready (cmpi29_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork90_outs_8, fork90_outs_7, fork90_outs_6, fork90_outs_5, fork90_outs_4, fork90_outs_3, fork90_outs_2, fork90_outs_1, fork90_outs_0}),
    .outs_valid ({fork90_outs_8_valid, fork90_outs_7_valid, fork90_outs_6_valid, fork90_outs_5_valid, fork90_outs_4_valid, fork90_outs_3_valid, fork90_outs_2_valid, fork90_outs_1_valid, fork90_outs_0_valid}),
    .outs_ready ({fork90_outs_8_ready, fork90_outs_7_ready, fork90_outs_6_ready, fork90_outs_5_ready, fork90_outs_4_ready, fork90_outs_3_ready, fork90_outs_2_ready, fork90_outs_1_ready, fork90_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br293(
    .condition (fork90_outs_4),
    .condition_valid (fork90_outs_4_valid),
    .condition_ready (fork90_outs_4_ready),
    .data (constant426_outs),
    .data_valid (constant426_outs_valid),
    .data_ready (constant426_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br293_trueOut),
    .trueOut_valid (cond_br293_trueOut_valid),
    .trueOut_ready (cond_br293_trueOut_ready),
    .falseOut (cond_br293_falseOut),
    .falseOut_valid (cond_br293_falseOut_valid),
    .falseOut_ready (cond_br293_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink232(
    .ins (cond_br293_falseOut),
    .ins_valid (cond_br293_falseOut_valid),
    .ins_ready (cond_br293_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br294(
    .condition (fork90_outs_7),
    .condition_valid (fork90_outs_7_valid),
    .condition_ready (fork90_outs_7_ready),
    .data (constant560_outs),
    .data_valid (constant560_outs_valid),
    .data_ready (constant560_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br294_trueOut),
    .trueOut_valid (cond_br294_trueOut_valid),
    .trueOut_ready (cond_br294_trueOut_ready),
    .falseOut (cond_br294_falseOut),
    .falseOut_valid (cond_br294_falseOut_valid),
    .falseOut_ready (cond_br294_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink233(
    .ins (cond_br294_falseOut),
    .ins_valid (cond_br294_falseOut_valid),
    .ins_ready (cond_br294_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(27), .OUTPUT_TYPE(33)) extsi234(
    .ins (cond_br294_trueOut),
    .ins_valid (cond_br294_trueOut_valid),
    .ins_ready (cond_br294_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi234_outs),
    .outs_valid (extsi234_outs_valid),
    .outs_ready (extsi234_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br295(
    .condition (fork90_outs_3),
    .condition_valid (fork90_outs_3_valid),
    .condition_ready (fork90_outs_3_ready),
    .data (constant428_outs),
    .data_valid (constant428_outs_valid),
    .data_ready (constant428_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br295_trueOut),
    .trueOut_valid (cond_br295_trueOut_valid),
    .trueOut_ready (cond_br295_trueOut_ready),
    .falseOut (cond_br295_falseOut),
    .falseOut_valid (cond_br295_falseOut_valid),
    .falseOut_ready (cond_br295_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink234(
    .ins (cond_br295_falseOut),
    .ins_valid (cond_br295_falseOut_valid),
    .ins_ready (cond_br295_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(17)) cond_br296(
    .condition (fork90_outs_6),
    .condition_valid (fork90_outs_6_valid),
    .condition_ready (fork90_outs_6_ready),
    .data (constant561_outs),
    .data_valid (constant561_outs_valid),
    .data_ready (constant561_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br296_trueOut),
    .trueOut_valid (cond_br296_trueOut_valid),
    .trueOut_ready (cond_br296_trueOut_ready),
    .falseOut (cond_br296_falseOut),
    .falseOut_valid (cond_br296_falseOut_valid),
    .falseOut_ready (cond_br296_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink235(
    .ins (cond_br296_falseOut),
    .ins_valid (cond_br296_falseOut_valid),
    .ins_ready (cond_br296_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(17), .OUTPUT_TYPE(22)) extsi235(
    .ins (cond_br296_trueOut),
    .ins_valid (cond_br296_trueOut_valid),
    .ins_ready (cond_br296_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi235_outs),
    .outs_valid (extsi235_outs_valid),
    .outs_ready (extsi235_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br297(
    .condition (fork90_outs_2),
    .condition_valid (fork90_outs_2_valid),
    .condition_ready (fork90_outs_2_ready),
    .data (constant430_outs),
    .data_valid (constant430_outs_valid),
    .data_ready (constant430_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br297_trueOut),
    .trueOut_valid (cond_br297_trueOut_valid),
    .trueOut_ready (cond_br297_trueOut_ready),
    .falseOut (cond_br297_falseOut),
    .falseOut_valid (cond_br297_falseOut_valid),
    .falseOut_ready (cond_br297_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink236(
    .ins (cond_br297_falseOut),
    .ins_valid (cond_br297_falseOut_valid),
    .ins_ready (cond_br297_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(6)) cond_br298(
    .condition (fork90_outs_5),
    .condition_valid (fork90_outs_5_valid),
    .condition_ready (fork90_outs_5_ready),
    .data (constant562_outs),
    .data_valid (constant562_outs_valid),
    .data_ready (constant562_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br298_trueOut),
    .trueOut_valid (cond_br298_trueOut_valid),
    .trueOut_ready (cond_br298_trueOut_ready),
    .falseOut (cond_br298_falseOut),
    .falseOut_valid (cond_br298_falseOut_valid),
    .falseOut_ready (cond_br298_falseOut_ready)
  );

  sink #(.DATA_TYPE(6)) sink237(
    .ins (cond_br298_falseOut),
    .ins_valid (cond_br298_falseOut_valid),
    .ins_ready (cond_br298_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(12)) extsi236(
    .ins (cond_br298_trueOut),
    .ins_valid (cond_br298_trueOut_valid),
    .ins_ready (cond_br298_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi236_outs),
    .outs_valid (extsi236_outs_valid),
    .outs_ready (extsi236_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer168(
    .ins (cond_br290_falseOut),
    .ins_valid (cond_br290_falseOut_valid),
    .ins_ready (cond_br290_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer168_outs),
    .outs_valid (buffer168_outs_valid),
    .outs_ready (buffer168_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer169(
    .ins (buffer168_outs),
    .ins_valid (buffer168_outs_valid),
    .ins_ready (buffer168_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer169_outs),
    .outs_valid (buffer169_outs_valid),
    .outs_ready (buffer169_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br299(
    .condition (fork90_outs_0),
    .condition_valid (fork90_outs_0_valid),
    .condition_ready (fork90_outs_0_ready),
    .data (buffer169_outs),
    .data_valid (buffer169_outs_valid),
    .data_ready (buffer169_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br299_trueOut),
    .trueOut_valid (cond_br299_trueOut_valid),
    .trueOut_ready (cond_br299_trueOut_ready),
    .falseOut (cond_br299_falseOut),
    .falseOut_valid (cond_br299_falseOut_valid),
    .falseOut_ready (cond_br299_falseOut_ready)
  );

  cond_br_dataless cond_br300(
    .condition (fork90_outs_1),
    .condition_valid (fork90_outs_1_valid),
    .condition_ready (fork90_outs_1_ready),
    .data_valid (fork89_outs_6_valid),
    .data_ready (fork89_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br300_trueOut_valid),
    .trueOut_ready (cond_br300_trueOut_ready),
    .falseOut_valid (cond_br300_falseOut_valid),
    .falseOut_ready (cond_br300_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br301(
    .condition (fork90_outs_8),
    .condition_valid (fork90_outs_8_valid),
    .condition_ready (fork90_outs_8_ready),
    .data (fork88_outs_1),
    .data_valid (fork88_outs_1_valid),
    .data_ready (fork88_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br301_trueOut),
    .trueOut_valid (cond_br301_trueOut_valid),
    .trueOut_ready (cond_br301_trueOut_ready),
    .falseOut (cond_br301_falseOut),
    .falseOut_valid (cond_br301_falseOut_valid),
    .falseOut_ready (cond_br301_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink238(
    .ins (cond_br301_trueOut),
    .ins_valid (cond_br301_trueOut_valid),
    .ins_ready (cond_br301_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer176(
    .ins (cond_br301_falseOut),
    .ins_valid (cond_br301_falseOut_valid),
    .ins_ready (cond_br301_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer176_outs),
    .outs_valid (buffer176_outs_valid),
    .outs_ready (buffer176_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer177(
    .ins (buffer176_outs),
    .ins_valid (buffer176_outs_valid),
    .ins_ready (buffer176_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer177_outs),
    .outs_valid (buffer177_outs_valid),
    .outs_ready (buffer177_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(5)) fork91(
    .ins (buffer177_outs),
    .ins_valid (buffer177_outs_valid),
    .ins_ready (buffer177_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork91_outs_1, fork91_outs_0}),
    .outs_valid ({fork91_outs_1_valid, fork91_outs_0_valid}),
    .outs_ready ({fork91_outs_1_ready, fork91_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi237(
    .ins (fork91_outs_0),
    .ins_valid (fork91_outs_0_valid),
    .ins_ready (fork91_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi237_outs),
    .outs_valid (extsi237_outs_valid),
    .outs_ready (extsi237_outs_ready)
  );

  oehb_dataless buffer178(
    .ins_valid (cond_br300_falseOut_valid),
    .ins_ready (cond_br300_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer178_outs_valid),
    .outs_ready (buffer178_outs_ready)
  );

  tehb_dataless buffer179(
    .ins_valid (buffer178_outs_valid),
    .ins_ready (buffer178_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer179_outs_valid),
    .outs_ready (buffer179_outs_ready)
  );

  fork_dataless #(.SIZE(7)) fork92(
    .ins_valid (buffer179_outs_valid),
    .ins_ready (buffer179_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork92_outs_6_valid, fork92_outs_5_valid, fork92_outs_4_valid, fork92_outs_3_valid, fork92_outs_2_valid, fork92_outs_1_valid, fork92_outs_0_valid}),
    .outs_ready ({fork92_outs_6_ready, fork92_outs_5_ready, fork92_outs_4_ready, fork92_outs_3_ready, fork92_outs_2_ready, fork92_outs_1_ready, fork92_outs_0_ready})
  );

  handshake_constant_207 #(.DATA_WIDTH(37)) constant433(
    .ctrl_valid (fork92_outs_5_valid),
    .ctrl_ready (fork92_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant433_outs),
    .outs_valid (constant433_outs_valid),
    .outs_ready (constant433_outs_ready)
  );

  handshake_constant_208 #(.DATA_WIDTH(27)) constant564(
    .ctrl_valid (fork92_outs_2_valid),
    .ctrl_ready (fork92_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant564_outs),
    .outs_valid (constant564_outs_valid),
    .outs_ready (constant564_outs_ready)
  );

  handshake_constant_209 #(.DATA_WIDTH(27)) constant435(
    .ctrl_valid (fork92_outs_4_valid),
    .ctrl_ready (fork92_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant435_outs),
    .outs_valid (constant435_outs_valid),
    .outs_ready (constant435_outs_ready)
  );

  handshake_constant_210 #(.DATA_WIDTH(17)) constant565(
    .ctrl_valid (fork92_outs_1_valid),
    .ctrl_ready (fork92_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant565_outs),
    .outs_valid (constant565_outs_valid),
    .outs_ready (constant565_outs_ready)
  );

  handshake_constant_211 #(.DATA_WIDTH(17)) constant437(
    .ctrl_valid (fork92_outs_3_valid),
    .ctrl_ready (fork92_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant437_outs),
    .outs_valid (constant437_outs_valid),
    .outs_ready (constant437_outs_ready)
  );

  handshake_constant_173 #(.DATA_WIDTH(6)) constant566(
    .ctrl_valid (fork92_outs_0_valid),
    .ctrl_ready (fork92_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant566_outs),
    .outs_valid (constant566_outs_valid),
    .outs_ready (constant566_outs_ready)
  );

  source source31(
    .clk (clk),
    .rst (rst),
    .outs_valid (source31_outs_valid),
    .outs_ready (source31_outs_ready)
  );

  handshake_constant_212 #(.DATA_WIDTH(6)) constant567(
    .ctrl_valid (source31_outs_valid),
    .ctrl_ready (source31_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant567_outs),
    .outs_valid (constant567_outs_valid),
    .outs_ready (constant567_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi30(
    .lhs (extsi237_outs),
    .lhs_valid (extsi237_outs_valid),
    .lhs_ready (extsi237_outs_ready),
    .rhs (constant567_outs),
    .rhs_valid (constant567_outs_valid),
    .rhs_ready (constant567_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi30_result),
    .result_valid (cmpi30_result_valid),
    .result_ready (cmpi30_result_ready)
  );

  fork_type #(.SIZE(9), .DATA_TYPE(1)) fork93(
    .ins (cmpi30_result),
    .ins_valid (cmpi30_result_valid),
    .ins_ready (cmpi30_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork93_outs_8, fork93_outs_7, fork93_outs_6, fork93_outs_5, fork93_outs_4, fork93_outs_3, fork93_outs_2, fork93_outs_1, fork93_outs_0}),
    .outs_valid ({fork93_outs_8_valid, fork93_outs_7_valid, fork93_outs_6_valid, fork93_outs_5_valid, fork93_outs_4_valid, fork93_outs_3_valid, fork93_outs_2_valid, fork93_outs_1_valid, fork93_outs_0_valid}),
    .outs_ready ({fork93_outs_8_ready, fork93_outs_7_ready, fork93_outs_6_ready, fork93_outs_5_ready, fork93_outs_4_ready, fork93_outs_3_ready, fork93_outs_2_ready, fork93_outs_1_ready, fork93_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br302(
    .condition (fork93_outs_4),
    .condition_valid (fork93_outs_4_valid),
    .condition_ready (fork93_outs_4_ready),
    .data (constant433_outs),
    .data_valid (constant433_outs_valid),
    .data_ready (constant433_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br302_trueOut),
    .trueOut_valid (cond_br302_trueOut_valid),
    .trueOut_ready (cond_br302_trueOut_ready),
    .falseOut (cond_br302_falseOut),
    .falseOut_valid (cond_br302_falseOut_valid),
    .falseOut_ready (cond_br302_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink240(
    .ins (cond_br302_falseOut),
    .ins_valid (cond_br302_falseOut_valid),
    .ins_ready (cond_br302_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br303(
    .condition (fork93_outs_7),
    .condition_valid (fork93_outs_7_valid),
    .condition_ready (fork93_outs_7_ready),
    .data (constant564_outs),
    .data_valid (constant564_outs_valid),
    .data_ready (constant564_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br303_trueOut),
    .trueOut_valid (cond_br303_trueOut_valid),
    .trueOut_ready (cond_br303_trueOut_ready),
    .falseOut (cond_br303_falseOut),
    .falseOut_valid (cond_br303_falseOut_valid),
    .falseOut_ready (cond_br303_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink241(
    .ins (cond_br303_falseOut),
    .ins_valid (cond_br303_falseOut_valid),
    .ins_ready (cond_br303_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(27), .OUTPUT_TYPE(33)) extsi238(
    .ins (cond_br303_trueOut),
    .ins_valid (cond_br303_trueOut_valid),
    .ins_ready (cond_br303_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi238_outs),
    .outs_valid (extsi238_outs_valid),
    .outs_ready (extsi238_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br304(
    .condition (fork93_outs_3),
    .condition_valid (fork93_outs_3_valid),
    .condition_ready (fork93_outs_3_ready),
    .data (constant435_outs),
    .data_valid (constant435_outs_valid),
    .data_ready (constant435_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br304_trueOut),
    .trueOut_valid (cond_br304_trueOut_valid),
    .trueOut_ready (cond_br304_trueOut_ready),
    .falseOut (cond_br304_falseOut),
    .falseOut_valid (cond_br304_falseOut_valid),
    .falseOut_ready (cond_br304_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink242(
    .ins (cond_br304_falseOut),
    .ins_valid (cond_br304_falseOut_valid),
    .ins_ready (cond_br304_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(17)) cond_br305(
    .condition (fork93_outs_6),
    .condition_valid (fork93_outs_6_valid),
    .condition_ready (fork93_outs_6_ready),
    .data (constant565_outs),
    .data_valid (constant565_outs_valid),
    .data_ready (constant565_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br305_trueOut),
    .trueOut_valid (cond_br305_trueOut_valid),
    .trueOut_ready (cond_br305_trueOut_ready),
    .falseOut (cond_br305_falseOut),
    .falseOut_valid (cond_br305_falseOut_valid),
    .falseOut_ready (cond_br305_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink243(
    .ins (cond_br305_falseOut),
    .ins_valid (cond_br305_falseOut_valid),
    .ins_ready (cond_br305_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(17), .OUTPUT_TYPE(22)) extsi239(
    .ins (cond_br305_trueOut),
    .ins_valid (cond_br305_trueOut_valid),
    .ins_ready (cond_br305_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi239_outs),
    .outs_valid (extsi239_outs_valid),
    .outs_ready (extsi239_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br306(
    .condition (fork93_outs_2),
    .condition_valid (fork93_outs_2_valid),
    .condition_ready (fork93_outs_2_ready),
    .data (constant437_outs),
    .data_valid (constant437_outs_valid),
    .data_ready (constant437_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br306_trueOut),
    .trueOut_valid (cond_br306_trueOut_valid),
    .trueOut_ready (cond_br306_trueOut_ready),
    .falseOut (cond_br306_falseOut),
    .falseOut_valid (cond_br306_falseOut_valid),
    .falseOut_ready (cond_br306_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink244(
    .ins (cond_br306_falseOut),
    .ins_valid (cond_br306_falseOut_valid),
    .ins_ready (cond_br306_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(6)) cond_br307(
    .condition (fork93_outs_5),
    .condition_valid (fork93_outs_5_valid),
    .condition_ready (fork93_outs_5_ready),
    .data (constant566_outs),
    .data_valid (constant566_outs_valid),
    .data_ready (constant566_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br307_trueOut),
    .trueOut_valid (cond_br307_trueOut_valid),
    .trueOut_ready (cond_br307_trueOut_ready),
    .falseOut (cond_br307_falseOut),
    .falseOut_valid (cond_br307_falseOut_valid),
    .falseOut_ready (cond_br307_falseOut_ready)
  );

  sink #(.DATA_TYPE(6)) sink245(
    .ins (cond_br307_falseOut),
    .ins_valid (cond_br307_falseOut_valid),
    .ins_ready (cond_br307_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(12)) extsi240(
    .ins (cond_br307_trueOut),
    .ins_valid (cond_br307_trueOut_valid),
    .ins_ready (cond_br307_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi240_outs),
    .outs_valid (extsi240_outs_valid),
    .outs_ready (extsi240_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer174(
    .ins (cond_br299_falseOut),
    .ins_valid (cond_br299_falseOut_valid),
    .ins_ready (cond_br299_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer174_outs),
    .outs_valid (buffer174_outs_valid),
    .outs_ready (buffer174_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer175(
    .ins (buffer174_outs),
    .ins_valid (buffer174_outs_valid),
    .ins_ready (buffer174_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer175_outs),
    .outs_valid (buffer175_outs_valid),
    .outs_ready (buffer175_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br308(
    .condition (fork93_outs_0),
    .condition_valid (fork93_outs_0_valid),
    .condition_ready (fork93_outs_0_ready),
    .data (buffer175_outs),
    .data_valid (buffer175_outs_valid),
    .data_ready (buffer175_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br308_trueOut),
    .trueOut_valid (cond_br308_trueOut_valid),
    .trueOut_ready (cond_br308_trueOut_ready),
    .falseOut (cond_br308_falseOut),
    .falseOut_valid (cond_br308_falseOut_valid),
    .falseOut_ready (cond_br308_falseOut_ready)
  );

  cond_br_dataless cond_br309(
    .condition (fork93_outs_1),
    .condition_valid (fork93_outs_1_valid),
    .condition_ready (fork93_outs_1_ready),
    .data_valid (fork92_outs_6_valid),
    .data_ready (fork92_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br309_trueOut_valid),
    .trueOut_ready (cond_br309_trueOut_ready),
    .falseOut_valid (cond_br309_falseOut_valid),
    .falseOut_ready (cond_br309_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(5)) cond_br310(
    .condition (fork93_outs_8),
    .condition_valid (fork93_outs_8_valid),
    .condition_ready (fork93_outs_8_ready),
    .data (fork91_outs_1),
    .data_valid (fork91_outs_1_valid),
    .data_ready (fork91_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br310_trueOut),
    .trueOut_valid (cond_br310_trueOut_valid),
    .trueOut_ready (cond_br310_trueOut_ready),
    .falseOut (cond_br310_falseOut),
    .falseOut_valid (cond_br310_falseOut_valid),
    .falseOut_ready (cond_br310_falseOut_ready)
  );

  sink #(.DATA_TYPE(5)) sink246(
    .ins (cond_br310_trueOut),
    .ins_valid (cond_br310_trueOut_valid),
    .ins_ready (cond_br310_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(5)) buffer182(
    .ins (cond_br310_falseOut),
    .ins_valid (cond_br310_falseOut_valid),
    .ins_ready (cond_br310_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer182_outs),
    .outs_valid (buffer182_outs_valid),
    .outs_ready (buffer182_outs_ready)
  );

  tehb #(.DATA_TYPE(5)) buffer183(
    .ins (buffer182_outs),
    .ins_valid (buffer182_outs_valid),
    .ins_ready (buffer182_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer183_outs),
    .outs_valid (buffer183_outs_valid),
    .outs_ready (buffer183_outs_ready)
  );

  extsi #(.INPUT_TYPE(5), .OUTPUT_TYPE(6)) extsi241(
    .ins (buffer183_outs),
    .ins_valid (buffer183_outs_valid),
    .ins_ready (buffer183_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi241_outs),
    .outs_valid (extsi241_outs_valid),
    .outs_ready (extsi241_outs_ready)
  );

  oehb_dataless buffer184(
    .ins_valid (cond_br309_falseOut_valid),
    .ins_ready (cond_br309_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer184_outs_valid),
    .outs_ready (buffer184_outs_ready)
  );

  tehb_dataless buffer185(
    .ins_valid (buffer184_outs_valid),
    .ins_ready (buffer184_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer185_outs_valid),
    .outs_ready (buffer185_outs_ready)
  );

  fork_dataless #(.SIZE(13)) fork94(
    .ins_valid (buffer185_outs_valid),
    .ins_ready (buffer185_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork94_outs_12_valid, fork94_outs_11_valid, fork94_outs_10_valid, fork94_outs_9_valid, fork94_outs_8_valid, fork94_outs_7_valid, fork94_outs_6_valid, fork94_outs_5_valid, fork94_outs_4_valid, fork94_outs_3_valid, fork94_outs_2_valid, fork94_outs_1_valid, fork94_outs_0_valid}),
    .outs_ready ({fork94_outs_12_ready, fork94_outs_11_ready, fork94_outs_10_ready, fork94_outs_9_ready, fork94_outs_8_ready, fork94_outs_7_ready, fork94_outs_6_ready, fork94_outs_5_ready, fork94_outs_4_ready, fork94_outs_3_ready, fork94_outs_2_ready, fork94_outs_1_ready, fork94_outs_0_ready})
  );

  handshake_constant_6 #(.DATA_WIDTH(33)) constant568(
    .ctrl_valid (fork94_outs_4_valid),
    .ctrl_ready (fork94_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant568_outs),
    .outs_valid (constant568_outs_valid),
    .outs_ready (constant568_outs_ready)
  );

  handshake_constant_5 #(.DATA_WIDTH(33)) constant441(
    .ctrl_valid (fork94_outs_11_valid),
    .ctrl_ready (fork94_outs_11_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant441_outs),
    .outs_valid (constant441_outs_valid),
    .outs_ready (constant441_outs_ready)
  );

  handshake_constant_4 #(.DATA_WIDTH(27)) constant442(
    .ctrl_valid (fork94_outs_10_valid),
    .ctrl_ready (fork94_outs_10_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant442_outs),
    .outs_valid (constant442_outs_valid),
    .outs_ready (constant442_outs_ready)
  );

  handshake_constant_3 #(.DATA_WIDTH(22)) constant443(
    .ctrl_valid (fork94_outs_9_valid),
    .ctrl_ready (fork94_outs_9_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant443_outs),
    .outs_valid (constant443_outs_valid),
    .outs_ready (constant443_outs_ready)
  );

  handshake_constant_2 #(.DATA_WIDTH(15)) constant569(
    .ctrl_valid (fork94_outs_3_valid),
    .ctrl_ready (fork94_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant569_outs),
    .outs_valid (constant569_outs_valid),
    .outs_ready (constant569_outs_ready)
  );

  handshake_constant_1 #(.DATA_WIDTH(12)) constant445(
    .ctrl_valid (fork94_outs_8_valid),
    .ctrl_ready (fork94_outs_8_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant445_outs),
    .outs_valid (constant445_outs_valid),
    .outs_ready (constant445_outs_ready)
  );

  handshake_constant_213 #(.DATA_WIDTH(37)) constant446(
    .ctrl_valid (fork94_outs_7_valid),
    .ctrl_ready (fork94_outs_7_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant446_outs),
    .outs_valid (constant446_outs_valid),
    .outs_ready (constant446_outs_ready)
  );

  handshake_constant_214 #(.DATA_WIDTH(26)) constant570(
    .ctrl_valid (fork94_outs_2_valid),
    .ctrl_ready (fork94_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant570_outs),
    .outs_valid (constant570_outs_valid),
    .outs_ready (constant570_outs_ready)
  );

  handshake_constant_215 #(.DATA_WIDTH(27)) constant448(
    .ctrl_valid (fork94_outs_6_valid),
    .ctrl_ready (fork94_outs_6_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant448_outs),
    .outs_valid (constant448_outs_valid),
    .outs_ready (constant448_outs_ready)
  );

  handshake_constant_216 #(.DATA_WIDTH(17)) constant571(
    .ctrl_valid (fork94_outs_1_valid),
    .ctrl_ready (fork94_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant571_outs),
    .outs_valid (constant571_outs_valid),
    .outs_ready (constant571_outs_ready)
  );

  handshake_constant_217 #(.DATA_WIDTH(17)) constant450(
    .ctrl_valid (fork94_outs_5_valid),
    .ctrl_ready (fork94_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant450_outs),
    .outs_valid (constant450_outs_valid),
    .outs_ready (constant450_outs_ready)
  );

  handshake_constant_146 #(.DATA_WIDTH(6)) constant572(
    .ctrl_valid (fork94_outs_0_valid),
    .ctrl_ready (fork94_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant572_outs),
    .outs_valid (constant572_outs_valid),
    .outs_ready (constant572_outs_ready)
  );

  source source32(
    .clk (clk),
    .rst (rst),
    .outs_valid (source32_outs_valid),
    .outs_ready (source32_outs_ready)
  );

  handshake_constant_199 #(.DATA_WIDTH(6)) constant573(
    .ctrl_valid (source32_outs_valid),
    .ctrl_ready (source32_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant573_outs),
    .outs_valid (constant573_outs_valid),
    .outs_ready (constant573_outs_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(6)) cmpi31(
    .lhs (extsi241_outs),
    .lhs_valid (extsi241_outs_valid),
    .lhs_ready (extsi241_outs_ready),
    .rhs (constant573_outs),
    .rhs_valid (constant573_outs_valid),
    .rhs_ready (constant573_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi31_result),
    .result_valid (cmpi31_result_valid),
    .result_ready (cmpi31_result_ready)
  );

  fork_type #(.SIZE(14), .DATA_TYPE(1)) fork95(
    .ins (cmpi31_result),
    .ins_valid (cmpi31_result_valid),
    .ins_ready (cmpi31_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork95_outs_13, fork95_outs_12, fork95_outs_11, fork95_outs_10, fork95_outs_9, fork95_outs_8, fork95_outs_7, fork95_outs_6, fork95_outs_5, fork95_outs_4, fork95_outs_3, fork95_outs_2, fork95_outs_1, fork95_outs_0}),
    .outs_valid ({fork95_outs_13_valid, fork95_outs_12_valid, fork95_outs_11_valid, fork95_outs_10_valid, fork95_outs_9_valid, fork95_outs_8_valid, fork95_outs_7_valid, fork95_outs_6_valid, fork95_outs_5_valid, fork95_outs_4_valid, fork95_outs_3_valid, fork95_outs_2_valid, fork95_outs_1_valid, fork95_outs_0_valid}),
    .outs_ready ({fork95_outs_13_ready, fork95_outs_12_ready, fork95_outs_11_ready, fork95_outs_10_ready, fork95_outs_9_ready, fork95_outs_8_ready, fork95_outs_7_ready, fork95_outs_6_ready, fork95_outs_5_ready, fork95_outs_4_ready, fork95_outs_3_ready, fork95_outs_2_ready, fork95_outs_1_ready, fork95_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(37)) cond_br311(
    .condition (fork95_outs_8),
    .condition_valid (fork95_outs_8_valid),
    .condition_ready (fork95_outs_8_ready),
    .data (constant446_outs),
    .data_valid (constant446_outs_valid),
    .data_ready (constant446_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br311_trueOut),
    .trueOut_valid (cond_br311_trueOut_valid),
    .trueOut_ready (cond_br311_trueOut_ready),
    .falseOut (cond_br311_falseOut),
    .falseOut_valid (cond_br311_falseOut_valid),
    .falseOut_ready (cond_br311_falseOut_ready)
  );

  sink #(.DATA_TYPE(37)) sink248(
    .ins (cond_br311_falseOut),
    .ins_valid (cond_br311_falseOut_valid),
    .ins_ready (cond_br311_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(26)) cond_br312(
    .condition (fork95_outs_13),
    .condition_valid (fork95_outs_13_valid),
    .condition_ready (fork95_outs_13_ready),
    .data (constant570_outs),
    .data_valid (constant570_outs_valid),
    .data_ready (constant570_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br312_trueOut),
    .trueOut_valid (cond_br312_trueOut_valid),
    .trueOut_ready (cond_br312_trueOut_ready),
    .falseOut (cond_br312_falseOut),
    .falseOut_valid (cond_br312_falseOut_valid),
    .falseOut_ready (cond_br312_falseOut_ready)
  );

  sink #(.DATA_TYPE(26)) sink249(
    .ins (cond_br312_falseOut),
    .ins_valid (cond_br312_falseOut_valid),
    .ins_ready (cond_br312_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(26), .OUTPUT_TYPE(33)) extsi242(
    .ins (cond_br312_trueOut),
    .ins_valid (cond_br312_trueOut_valid),
    .ins_ready (cond_br312_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi242_outs),
    .outs_valid (extsi242_outs_valid),
    .outs_ready (extsi242_outs_ready)
  );

  cond_br #(.DATA_TYPE(27)) cond_br313(
    .condition (fork95_outs_7),
    .condition_valid (fork95_outs_7_valid),
    .condition_ready (fork95_outs_7_ready),
    .data (constant448_outs),
    .data_valid (constant448_outs_valid),
    .data_ready (constant448_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br313_trueOut),
    .trueOut_valid (cond_br313_trueOut_valid),
    .trueOut_ready (cond_br313_trueOut_ready),
    .falseOut (cond_br313_falseOut),
    .falseOut_valid (cond_br313_falseOut_valid),
    .falseOut_ready (cond_br313_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink250(
    .ins (cond_br313_falseOut),
    .ins_valid (cond_br313_falseOut_valid),
    .ins_ready (cond_br313_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(17)) cond_br314(
    .condition (fork95_outs_12),
    .condition_valid (fork95_outs_12_valid),
    .condition_ready (fork95_outs_12_ready),
    .data (constant571_outs),
    .data_valid (constant571_outs_valid),
    .data_ready (constant571_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br314_trueOut),
    .trueOut_valid (cond_br314_trueOut_valid),
    .trueOut_ready (cond_br314_trueOut_ready),
    .falseOut (cond_br314_falseOut),
    .falseOut_valid (cond_br314_falseOut_valid),
    .falseOut_ready (cond_br314_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink251(
    .ins (cond_br314_falseOut),
    .ins_valid (cond_br314_falseOut_valid),
    .ins_ready (cond_br314_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(17), .OUTPUT_TYPE(22)) extsi243(
    .ins (cond_br314_trueOut),
    .ins_valid (cond_br314_trueOut_valid),
    .ins_ready (cond_br314_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi243_outs),
    .outs_valid (extsi243_outs_valid),
    .outs_ready (extsi243_outs_ready)
  );

  cond_br #(.DATA_TYPE(17)) cond_br315(
    .condition (fork95_outs_6),
    .condition_valid (fork95_outs_6_valid),
    .condition_ready (fork95_outs_6_ready),
    .data (constant450_outs),
    .data_valid (constant450_outs_valid),
    .data_ready (constant450_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br315_trueOut),
    .trueOut_valid (cond_br315_trueOut_valid),
    .trueOut_ready (cond_br315_trueOut_ready),
    .falseOut (cond_br315_falseOut),
    .falseOut_valid (cond_br315_falseOut_valid),
    .falseOut_ready (cond_br315_falseOut_ready)
  );

  sink #(.DATA_TYPE(17)) sink252(
    .ins (cond_br315_falseOut),
    .ins_valid (cond_br315_falseOut_valid),
    .ins_ready (cond_br315_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(6)) cond_br316(
    .condition (fork95_outs_11),
    .condition_valid (fork95_outs_11_valid),
    .condition_ready (fork95_outs_11_ready),
    .data (constant572_outs),
    .data_valid (constant572_outs_valid),
    .data_ready (constant572_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br316_trueOut),
    .trueOut_valid (cond_br316_trueOut_valid),
    .trueOut_ready (cond_br316_trueOut_ready),
    .falseOut (cond_br316_falseOut),
    .falseOut_valid (cond_br316_falseOut_valid),
    .falseOut_ready (cond_br316_falseOut_ready)
  );

  sink #(.DATA_TYPE(6)) sink253(
    .ins (cond_br316_falseOut),
    .ins_valid (cond_br316_falseOut_valid),
    .ins_ready (cond_br316_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(12)) extsi244(
    .ins (cond_br316_trueOut),
    .ins_valid (cond_br316_trueOut_valid),
    .ins_ready (cond_br316_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi244_outs),
    .outs_valid (extsi244_outs_valid),
    .outs_ready (extsi244_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer180(
    .ins (cond_br308_falseOut),
    .ins_valid (cond_br308_falseOut_valid),
    .ins_ready (cond_br308_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer180_outs),
    .outs_valid (buffer180_outs_valid),
    .outs_ready (buffer180_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer181(
    .ins (buffer180_outs),
    .ins_valid (buffer180_outs_valid),
    .ins_ready (buffer180_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer181_outs),
    .outs_valid (buffer181_outs_valid),
    .outs_ready (buffer181_outs_ready)
  );

  cond_br #(.DATA_TYPE(7)) cond_br317(
    .condition (fork95_outs_0),
    .condition_valid (fork95_outs_0_valid),
    .condition_ready (fork95_outs_0_ready),
    .data (buffer181_outs),
    .data_valid (buffer181_outs_valid),
    .data_ready (buffer181_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br317_trueOut),
    .trueOut_valid (cond_br317_trueOut_valid),
    .trueOut_ready (cond_br317_trueOut_ready),
    .falseOut (cond_br317_falseOut),
    .falseOut_valid (cond_br317_falseOut_valid),
    .falseOut_ready (cond_br317_falseOut_ready)
  );

  sink #(.DATA_TYPE(7)) sink254(
    .ins (cond_br317_falseOut),
    .ins_valid (cond_br317_falseOut_valid),
    .ins_ready (cond_br317_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(7)) fork96(
    .ins (cond_br317_trueOut),
    .ins_valid (cond_br317_trueOut_valid),
    .ins_ready (cond_br317_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork96_outs_1, fork96_outs_0}),
    .outs_valid ({fork96_outs_1_valid, fork96_outs_0_valid}),
    .outs_ready ({fork96_outs_1_ready, fork96_outs_0_ready})
  );

  cond_br_dataless cond_br318(
    .condition (fork95_outs_5),
    .condition_valid (fork95_outs_5_valid),
    .condition_ready (fork95_outs_5_ready),
    .data_valid (fork94_outs_12_valid),
    .data_ready (fork94_outs_12_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br318_trueOut_valid),
    .trueOut_ready (cond_br318_trueOut_ready),
    .falseOut_valid (cond_br318_falseOut_valid),
    .falseOut_ready (cond_br318_falseOut_ready)
  );

  sink_dataless sink255(
    .ins_valid (cond_br318_falseOut_valid),
    .ins_ready (cond_br318_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  fork_dataless #(.SIZE(2)) fork97(
    .ins_valid (cond_br318_trueOut_valid),
    .ins_ready (cond_br318_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork97_outs_1_valid, fork97_outs_0_valid}),
    .outs_ready ({fork97_outs_1_ready, fork97_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(33)) cond_br319(
    .condition (fork95_outs_10),
    .condition_valid (fork95_outs_10_valid),
    .condition_ready (fork95_outs_10_ready),
    .data (constant568_outs),
    .data_valid (constant568_outs_valid),
    .data_ready (constant568_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br319_trueOut),
    .trueOut_valid (cond_br319_trueOut_valid),
    .trueOut_ready (cond_br319_trueOut_ready),
    .falseOut (cond_br319_falseOut),
    .falseOut_valid (cond_br319_falseOut_valid),
    .falseOut_ready (cond_br319_falseOut_ready)
  );

  sink #(.DATA_TYPE(33)) sink256(
    .ins (cond_br319_falseOut),
    .ins_valid (cond_br319_falseOut_valid),
    .ins_ready (cond_br319_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(33), .OUTPUT_TYPE(37)) extsi245(
    .ins (cond_br319_trueOut),
    .ins_valid (cond_br319_trueOut_valid),
    .ins_ready (cond_br319_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi245_outs),
    .outs_valid (extsi245_outs_valid),
    .outs_ready (extsi245_outs_ready)
  );

  cond_br #(.DATA_TYPE(33)) cond_br320(
    .condition (fork95_outs_4),
    .condition_valid (fork95_outs_4_valid),
    .condition_ready (fork95_outs_4_ready),
    .data (constant441_outs),
    .data_valid (constant441_outs_valid),
    .data_ready (constant441_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br320_trueOut),
    .trueOut_valid (cond_br320_trueOut_valid),
    .trueOut_ready (cond_br320_trueOut_ready),
    .falseOut (cond_br320_falseOut),
    .falseOut_valid (cond_br320_falseOut_valid),
    .falseOut_ready (cond_br320_falseOut_ready)
  );

  sink #(.DATA_TYPE(33)) sink257(
    .ins (cond_br320_falseOut),
    .ins_valid (cond_br320_falseOut_valid),
    .ins_ready (cond_br320_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(27)) cond_br321(
    .condition (fork95_outs_3),
    .condition_valid (fork95_outs_3_valid),
    .condition_ready (fork95_outs_3_ready),
    .data (constant442_outs),
    .data_valid (constant442_outs_valid),
    .data_ready (constant442_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br321_trueOut),
    .trueOut_valid (cond_br321_trueOut_valid),
    .trueOut_ready (cond_br321_trueOut_ready),
    .falseOut (cond_br321_falseOut),
    .falseOut_valid (cond_br321_falseOut_valid),
    .falseOut_ready (cond_br321_falseOut_ready)
  );

  sink #(.DATA_TYPE(27)) sink258(
    .ins (cond_br321_falseOut),
    .ins_valid (cond_br321_falseOut_valid),
    .ins_ready (cond_br321_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(22)) cond_br322(
    .condition (fork95_outs_2),
    .condition_valid (fork95_outs_2_valid),
    .condition_ready (fork95_outs_2_ready),
    .data (constant443_outs),
    .data_valid (constant443_outs_valid),
    .data_ready (constant443_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br322_trueOut),
    .trueOut_valid (cond_br322_trueOut_valid),
    .trueOut_ready (cond_br322_trueOut_ready),
    .falseOut (cond_br322_falseOut),
    .falseOut_valid (cond_br322_falseOut_valid),
    .falseOut_ready (cond_br322_falseOut_ready)
  );

  sink #(.DATA_TYPE(22)) sink259(
    .ins (cond_br322_falseOut),
    .ins_valid (cond_br322_falseOut_valid),
    .ins_ready (cond_br322_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(15)) cond_br323(
    .condition (fork95_outs_9),
    .condition_valid (fork95_outs_9_valid),
    .condition_ready (fork95_outs_9_ready),
    .data (constant569_outs),
    .data_valid (constant569_outs_valid),
    .data_ready (constant569_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br323_trueOut),
    .trueOut_valid (cond_br323_trueOut_valid),
    .trueOut_ready (cond_br323_trueOut_ready),
    .falseOut (cond_br323_falseOut),
    .falseOut_valid (cond_br323_falseOut_valid),
    .falseOut_ready (cond_br323_falseOut_ready)
  );

  sink #(.DATA_TYPE(15)) sink260(
    .ins (cond_br323_falseOut),
    .ins_valid (cond_br323_falseOut_valid),
    .ins_ready (cond_br323_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  extsi #(.INPUT_TYPE(15), .OUTPUT_TYPE(17)) extsi246(
    .ins (cond_br323_trueOut),
    .ins_valid (cond_br323_trueOut_valid),
    .ins_ready (cond_br323_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi246_outs),
    .outs_valid (extsi246_outs_valid),
    .outs_ready (extsi246_outs_ready)
  );

  cond_br #(.DATA_TYPE(12)) cond_br324(
    .condition (fork95_outs_1),
    .condition_valid (fork95_outs_1_valid),
    .condition_ready (fork95_outs_1_ready),
    .data (constant445_outs),
    .data_valid (constant445_outs_valid),
    .data_ready (constant445_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br324_trueOut),
    .trueOut_valid (cond_br324_trueOut_valid),
    .trueOut_ready (cond_br324_trueOut_ready),
    .falseOut (cond_br324_falseOut),
    .falseOut_valid (cond_br324_falseOut_valid),
    .falseOut_ready (cond_br324_falseOut_ready)
  );

  sink #(.DATA_TYPE(12)) sink261(
    .ins (cond_br324_falseOut),
    .ins_valid (cond_br324_falseOut_valid),
    .ins_ready (cond_br324_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  mux #(.SIZE(33), .DATA_TYPE(37), .SELECT_TYPE(6)) mux0(
    .index (fork99_outs_6),
    .index_valid (fork99_outs_6_valid),
    .index_ready (fork99_outs_6_ready),
    .ins ({extsi245_outs, cond_br311_trueOut, cond_br302_trueOut, cond_br293_trueOut, cond_br284_trueOut, cond_br275_trueOut, cond_br266_trueOut, cond_br257_trueOut, cond_br248_trueOut, cond_br239_trueOut, cond_br230_trueOut, cond_br221_trueOut, cond_br212_trueOut, cond_br203_trueOut, cond_br194_trueOut, cond_br185_trueOut, cond_br176_trueOut, cond_br167_trueOut, cond_br158_trueOut, cond_br149_trueOut, cond_br140_trueOut, cond_br131_trueOut, cond_br122_trueOut, cond_br113_trueOut, cond_br104_trueOut, cond_br95_trueOut, extsi157_outs, extsi155_outs, extsi153_outs, extsi150_outs, extsi148_outs, extsi145_outs, extsi142_outs}),
    .ins_valid ({extsi245_outs_valid, cond_br311_trueOut_valid, cond_br302_trueOut_valid, cond_br293_trueOut_valid, cond_br284_trueOut_valid, cond_br275_trueOut_valid, cond_br266_trueOut_valid, cond_br257_trueOut_valid, cond_br248_trueOut_valid, cond_br239_trueOut_valid, cond_br230_trueOut_valid, cond_br221_trueOut_valid, cond_br212_trueOut_valid, cond_br203_trueOut_valid, cond_br194_trueOut_valid, cond_br185_trueOut_valid, cond_br176_trueOut_valid, cond_br167_trueOut_valid, cond_br158_trueOut_valid, cond_br149_trueOut_valid, cond_br140_trueOut_valid, cond_br131_trueOut_valid, cond_br122_trueOut_valid, cond_br113_trueOut_valid, cond_br104_trueOut_valid, cond_br95_trueOut_valid, extsi157_outs_valid, extsi155_outs_valid, extsi153_outs_valid, extsi150_outs_valid, extsi148_outs_valid, extsi145_outs_valid, extsi142_outs_valid}),
    .ins_ready ({extsi245_outs_ready, cond_br311_trueOut_ready, cond_br302_trueOut_ready, cond_br293_trueOut_ready, cond_br284_trueOut_ready, cond_br275_trueOut_ready, cond_br266_trueOut_ready, cond_br257_trueOut_ready, cond_br248_trueOut_ready, cond_br239_trueOut_ready, cond_br230_trueOut_ready, cond_br221_trueOut_ready, cond_br212_trueOut_ready, cond_br203_trueOut_ready, cond_br194_trueOut_ready, cond_br185_trueOut_ready, cond_br176_trueOut_ready, cond_br167_trueOut_ready, cond_br158_trueOut_ready, cond_br149_trueOut_ready, cond_br140_trueOut_ready, cond_br131_trueOut_ready, cond_br122_trueOut_ready, cond_br113_trueOut_ready, cond_br104_trueOut_ready, cond_br95_trueOut_ready, extsi157_outs_ready, extsi155_outs_ready, extsi153_outs_ready, extsi150_outs_ready, extsi148_outs_ready, extsi145_outs_ready, extsi142_outs_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux0_outs),
    .outs_valid (mux0_outs_valid),
    .outs_ready (mux0_outs_ready)
  );

  mux #(.SIZE(33), .DATA_TYPE(33), .SELECT_TYPE(6)) mux1(
    .index (fork99_outs_5),
    .index_valid (fork99_outs_5_valid),
    .index_ready (fork99_outs_5_ready),
    .ins ({cond_br320_trueOut, extsi242_outs, extsi238_outs, extsi234_outs, extsi230_outs, extsi226_outs, extsi222_outs, extsi218_outs, extsi214_outs, extsi210_outs, extsi206_outs, extsi202_outs, extsi198_outs, extsi194_outs, extsi190_outs, extsi186_outs, extsi183_outs, extsi180_outs, extsi178_outs, extsi176_outs, extsi174_outs, extsi171_outs, extsi168_outs, extsi165_outs, extsi162_outs, extsi160_outs, extsi158_outs, cond_br78_trueOut, cond_br69_trueOut, cond_br60_trueOut, cond_br51_trueOut, cond_br42_trueOut, cond_br33_trueOut}),
    .ins_valid ({cond_br320_trueOut_valid, extsi242_outs_valid, extsi238_outs_valid, extsi234_outs_valid, extsi230_outs_valid, extsi226_outs_valid, extsi222_outs_valid, extsi218_outs_valid, extsi214_outs_valid, extsi210_outs_valid, extsi206_outs_valid, extsi202_outs_valid, extsi198_outs_valid, extsi194_outs_valid, extsi190_outs_valid, extsi186_outs_valid, extsi183_outs_valid, extsi180_outs_valid, extsi178_outs_valid, extsi176_outs_valid, extsi174_outs_valid, extsi171_outs_valid, extsi168_outs_valid, extsi165_outs_valid, extsi162_outs_valid, extsi160_outs_valid, extsi158_outs_valid, cond_br78_trueOut_valid, cond_br69_trueOut_valid, cond_br60_trueOut_valid, cond_br51_trueOut_valid, cond_br42_trueOut_valid, cond_br33_trueOut_valid}),
    .ins_ready ({cond_br320_trueOut_ready, extsi242_outs_ready, extsi238_outs_ready, extsi234_outs_ready, extsi230_outs_ready, extsi226_outs_ready, extsi222_outs_ready, extsi218_outs_ready, extsi214_outs_ready, extsi210_outs_ready, extsi206_outs_ready, extsi202_outs_ready, extsi198_outs_ready, extsi194_outs_ready, extsi190_outs_ready, extsi186_outs_ready, extsi183_outs_ready, extsi180_outs_ready, extsi178_outs_ready, extsi176_outs_ready, extsi174_outs_ready, extsi171_outs_ready, extsi168_outs_ready, extsi165_outs_ready, extsi162_outs_ready, extsi160_outs_ready, extsi158_outs_ready, cond_br78_trueOut_ready, cond_br69_trueOut_ready, cond_br60_trueOut_ready, cond_br51_trueOut_ready, cond_br42_trueOut_ready, cond_br33_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux1_outs),
    .outs_valid (mux1_outs_valid),
    .outs_ready (mux1_outs_ready)
  );

  mux #(.SIZE(33), .DATA_TYPE(27), .SELECT_TYPE(6)) mux2(
    .index (fork99_outs_4),
    .index_valid (fork99_outs_4_valid),
    .index_ready (fork99_outs_4_ready),
    .ins ({cond_br321_trueOut, cond_br313_trueOut, cond_br304_trueOut, cond_br295_trueOut, cond_br286_trueOut, cond_br277_trueOut, cond_br268_trueOut, cond_br259_trueOut, cond_br250_trueOut, cond_br241_trueOut, cond_br232_trueOut, cond_br223_trueOut, cond_br214_trueOut, cond_br205_trueOut, cond_br196_trueOut, cond_br187_trueOut, cond_br178_trueOut, cond_br169_trueOut, cond_br160_trueOut, cond_br151_trueOut, cond_br142_trueOut, cond_br133_trueOut, cond_br124_trueOut, cond_br115_trueOut, cond_br106_trueOut, cond_br97_trueOut, cond_br88_trueOut, cond_br79_trueOut, cond_br70_trueOut, cond_br61_trueOut, cond_br52_trueOut, cond_br43_trueOut, cond_br34_trueOut}),
    .ins_valid ({cond_br321_trueOut_valid, cond_br313_trueOut_valid, cond_br304_trueOut_valid, cond_br295_trueOut_valid, cond_br286_trueOut_valid, cond_br277_trueOut_valid, cond_br268_trueOut_valid, cond_br259_trueOut_valid, cond_br250_trueOut_valid, cond_br241_trueOut_valid, cond_br232_trueOut_valid, cond_br223_trueOut_valid, cond_br214_trueOut_valid, cond_br205_trueOut_valid, cond_br196_trueOut_valid, cond_br187_trueOut_valid, cond_br178_trueOut_valid, cond_br169_trueOut_valid, cond_br160_trueOut_valid, cond_br151_trueOut_valid, cond_br142_trueOut_valid, cond_br133_trueOut_valid, cond_br124_trueOut_valid, cond_br115_trueOut_valid, cond_br106_trueOut_valid, cond_br97_trueOut_valid, cond_br88_trueOut_valid, cond_br79_trueOut_valid, cond_br70_trueOut_valid, cond_br61_trueOut_valid, cond_br52_trueOut_valid, cond_br43_trueOut_valid, cond_br34_trueOut_valid}),
    .ins_ready ({cond_br321_trueOut_ready, cond_br313_trueOut_ready, cond_br304_trueOut_ready, cond_br295_trueOut_ready, cond_br286_trueOut_ready, cond_br277_trueOut_ready, cond_br268_trueOut_ready, cond_br259_trueOut_ready, cond_br250_trueOut_ready, cond_br241_trueOut_ready, cond_br232_trueOut_ready, cond_br223_trueOut_ready, cond_br214_trueOut_ready, cond_br205_trueOut_ready, cond_br196_trueOut_ready, cond_br187_trueOut_ready, cond_br178_trueOut_ready, cond_br169_trueOut_ready, cond_br160_trueOut_ready, cond_br151_trueOut_ready, cond_br142_trueOut_ready, cond_br133_trueOut_ready, cond_br124_trueOut_ready, cond_br115_trueOut_ready, cond_br106_trueOut_ready, cond_br97_trueOut_ready, cond_br88_trueOut_ready, cond_br79_trueOut_ready, cond_br70_trueOut_ready, cond_br61_trueOut_ready, cond_br52_trueOut_ready, cond_br43_trueOut_ready, cond_br34_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux2_outs),
    .outs_valid (mux2_outs_valid),
    .outs_ready (mux2_outs_ready)
  );

  mux #(.SIZE(33), .DATA_TYPE(22), .SELECT_TYPE(6)) mux3(
    .index (fork99_outs_3),
    .index_valid (fork99_outs_3_valid),
    .index_ready (fork99_outs_3_ready),
    .ins ({cond_br322_trueOut, extsi243_outs, extsi239_outs, extsi235_outs, extsi231_outs, extsi227_outs, extsi223_outs, extsi219_outs, extsi215_outs, extsi211_outs, extsi207_outs, extsi203_outs, extsi199_outs, extsi195_outs, extsi191_outs, extsi187_outs, extsi184_outs, extsi181_outs, extsi179_outs, extsi177_outs, extsi175_outs, extsi172_outs, extsi169_outs, extsi166_outs, extsi163_outs, extsi161_outs, cond_br89_trueOut, cond_br80_trueOut, cond_br71_trueOut, cond_br62_trueOut, cond_br53_trueOut, cond_br44_trueOut, cond_br35_trueOut}),
    .ins_valid ({cond_br322_trueOut_valid, extsi243_outs_valid, extsi239_outs_valid, extsi235_outs_valid, extsi231_outs_valid, extsi227_outs_valid, extsi223_outs_valid, extsi219_outs_valid, extsi215_outs_valid, extsi211_outs_valid, extsi207_outs_valid, extsi203_outs_valid, extsi199_outs_valid, extsi195_outs_valid, extsi191_outs_valid, extsi187_outs_valid, extsi184_outs_valid, extsi181_outs_valid, extsi179_outs_valid, extsi177_outs_valid, extsi175_outs_valid, extsi172_outs_valid, extsi169_outs_valid, extsi166_outs_valid, extsi163_outs_valid, extsi161_outs_valid, cond_br89_trueOut_valid, cond_br80_trueOut_valid, cond_br71_trueOut_valid, cond_br62_trueOut_valid, cond_br53_trueOut_valid, cond_br44_trueOut_valid, cond_br35_trueOut_valid}),
    .ins_ready ({cond_br322_trueOut_ready, extsi243_outs_ready, extsi239_outs_ready, extsi235_outs_ready, extsi231_outs_ready, extsi227_outs_ready, extsi223_outs_ready, extsi219_outs_ready, extsi215_outs_ready, extsi211_outs_ready, extsi207_outs_ready, extsi203_outs_ready, extsi199_outs_ready, extsi195_outs_ready, extsi191_outs_ready, extsi187_outs_ready, extsi184_outs_ready, extsi181_outs_ready, extsi179_outs_ready, extsi177_outs_ready, extsi175_outs_ready, extsi172_outs_ready, extsi169_outs_ready, extsi166_outs_ready, extsi163_outs_ready, extsi161_outs_ready, cond_br89_trueOut_ready, cond_br80_trueOut_ready, cond_br71_trueOut_ready, cond_br62_trueOut_ready, cond_br53_trueOut_ready, cond_br44_trueOut_ready, cond_br35_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux3_outs),
    .outs_valid (mux3_outs_valid),
    .outs_ready (mux3_outs_ready)
  );

  mux #(.SIZE(33), .DATA_TYPE(17), .SELECT_TYPE(6)) mux4(
    .index (fork99_outs_2),
    .index_valid (fork99_outs_2_valid),
    .index_ready (fork99_outs_2_ready),
    .ins ({extsi246_outs, cond_br315_trueOut, cond_br306_trueOut, cond_br297_trueOut, cond_br288_trueOut, cond_br279_trueOut, cond_br270_trueOut, cond_br261_trueOut, cond_br252_trueOut, cond_br243_trueOut, cond_br234_trueOut, cond_br225_trueOut, cond_br216_trueOut, cond_br207_trueOut, cond_br198_trueOut, cond_br189_trueOut, cond_br180_trueOut, cond_br171_trueOut, cond_br162_trueOut, cond_br153_trueOut, cond_br144_trueOut, extsi173_outs, extsi170_outs, extsi167_outs, extsi164_outs, cond_br99_trueOut, cond_br90_trueOut, cond_br81_trueOut, cond_br72_trueOut, cond_br63_trueOut, cond_br54_trueOut, extsi146_outs, extsi143_outs}),
    .ins_valid ({extsi246_outs_valid, cond_br315_trueOut_valid, cond_br306_trueOut_valid, cond_br297_trueOut_valid, cond_br288_trueOut_valid, cond_br279_trueOut_valid, cond_br270_trueOut_valid, cond_br261_trueOut_valid, cond_br252_trueOut_valid, cond_br243_trueOut_valid, cond_br234_trueOut_valid, cond_br225_trueOut_valid, cond_br216_trueOut_valid, cond_br207_trueOut_valid, cond_br198_trueOut_valid, cond_br189_trueOut_valid, cond_br180_trueOut_valid, cond_br171_trueOut_valid, cond_br162_trueOut_valid, cond_br153_trueOut_valid, cond_br144_trueOut_valid, extsi173_outs_valid, extsi170_outs_valid, extsi167_outs_valid, extsi164_outs_valid, cond_br99_trueOut_valid, cond_br90_trueOut_valid, cond_br81_trueOut_valid, cond_br72_trueOut_valid, cond_br63_trueOut_valid, cond_br54_trueOut_valid, extsi146_outs_valid, extsi143_outs_valid}),
    .ins_ready ({extsi246_outs_ready, cond_br315_trueOut_ready, cond_br306_trueOut_ready, cond_br297_trueOut_ready, cond_br288_trueOut_ready, cond_br279_trueOut_ready, cond_br270_trueOut_ready, cond_br261_trueOut_ready, cond_br252_trueOut_ready, cond_br243_trueOut_ready, cond_br234_trueOut_ready, cond_br225_trueOut_ready, cond_br216_trueOut_ready, cond_br207_trueOut_ready, cond_br198_trueOut_ready, cond_br189_trueOut_ready, cond_br180_trueOut_ready, cond_br171_trueOut_ready, cond_br162_trueOut_ready, cond_br153_trueOut_ready, cond_br144_trueOut_ready, extsi173_outs_ready, extsi170_outs_ready, extsi167_outs_ready, extsi164_outs_ready, cond_br99_trueOut_ready, cond_br90_trueOut_ready, cond_br81_trueOut_ready, cond_br72_trueOut_ready, cond_br63_trueOut_ready, cond_br54_trueOut_ready, extsi146_outs_ready, extsi143_outs_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux4_outs),
    .outs_valid (mux4_outs_valid),
    .outs_ready (mux4_outs_ready)
  );

  mux #(.SIZE(33), .DATA_TYPE(12), .SELECT_TYPE(6)) mux5(
    .index (fork99_outs_1),
    .index_valid (fork99_outs_1_valid),
    .index_ready (fork99_outs_1_ready),
    .ins ({cond_br324_trueOut, extsi244_outs, extsi240_outs, extsi236_outs, extsi232_outs, extsi228_outs, extsi224_outs, extsi220_outs, extsi216_outs, extsi212_outs, extsi208_outs, extsi204_outs, extsi200_outs, extsi196_outs, extsi192_outs, extsi188_outs, cond_br181_trueOut, cond_br172_trueOut, cond_br163_trueOut, cond_br154_trueOut, cond_br145_trueOut, cond_br136_trueOut, cond_br127_trueOut, cond_br118_trueOut, cond_br109_trueOut, cond_br100_trueOut, cond_br91_trueOut, cond_br82_trueOut, cond_br73_trueOut, extsi151_outs, cond_br55_trueOut, cond_br46_trueOut, cond_br37_trueOut}),
    .ins_valid ({cond_br324_trueOut_valid, extsi244_outs_valid, extsi240_outs_valid, extsi236_outs_valid, extsi232_outs_valid, extsi228_outs_valid, extsi224_outs_valid, extsi220_outs_valid, extsi216_outs_valid, extsi212_outs_valid, extsi208_outs_valid, extsi204_outs_valid, extsi200_outs_valid, extsi196_outs_valid, extsi192_outs_valid, extsi188_outs_valid, cond_br181_trueOut_valid, cond_br172_trueOut_valid, cond_br163_trueOut_valid, cond_br154_trueOut_valid, cond_br145_trueOut_valid, cond_br136_trueOut_valid, cond_br127_trueOut_valid, cond_br118_trueOut_valid, cond_br109_trueOut_valid, cond_br100_trueOut_valid, cond_br91_trueOut_valid, cond_br82_trueOut_valid, cond_br73_trueOut_valid, extsi151_outs_valid, cond_br55_trueOut_valid, cond_br46_trueOut_valid, cond_br37_trueOut_valid}),
    .ins_ready ({cond_br324_trueOut_ready, extsi244_outs_ready, extsi240_outs_ready, extsi236_outs_ready, extsi232_outs_ready, extsi228_outs_ready, extsi224_outs_ready, extsi220_outs_ready, extsi216_outs_ready, extsi212_outs_ready, extsi208_outs_ready, extsi204_outs_ready, extsi200_outs_ready, extsi196_outs_ready, extsi192_outs_ready, extsi188_outs_ready, cond_br181_trueOut_ready, cond_br172_trueOut_ready, cond_br163_trueOut_ready, cond_br154_trueOut_ready, cond_br145_trueOut_ready, cond_br136_trueOut_ready, cond_br127_trueOut_ready, cond_br118_trueOut_ready, cond_br109_trueOut_ready, cond_br100_trueOut_ready, cond_br91_trueOut_ready, cond_br82_trueOut_ready, cond_br73_trueOut_ready, extsi151_outs_ready, cond_br55_trueOut_ready, cond_br46_trueOut_ready, cond_br37_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux5_outs),
    .outs_valid (mux5_outs_valid),
    .outs_ready (mux5_outs_ready)
  );

  mux #(.SIZE(33), .DATA_TYPE(7), .SELECT_TYPE(6)) mux6(
    .index (fork99_outs_0),
    .index_valid (fork99_outs_0_valid),
    .index_ready (fork99_outs_0_ready),
    .ins ({fork96_outs_1, fork96_outs_0, cond_br308_trueOut, cond_br299_trueOut, cond_br290_trueOut, cond_br281_trueOut, cond_br272_trueOut, cond_br263_trueOut, cond_br254_trueOut, cond_br245_trueOut, cond_br236_trueOut, cond_br227_trueOut, cond_br218_trueOut, cond_br209_trueOut, cond_br200_trueOut, cond_br191_trueOut, cond_br182_trueOut, cond_br173_trueOut, cond_br164_trueOut, cond_br155_trueOut, cond_br146_trueOut, cond_br137_trueOut, cond_br128_trueOut, cond_br119_trueOut, cond_br110_trueOut, cond_br101_trueOut, cond_br92_trueOut, cond_br83_trueOut, cond_br74_trueOut, cond_br65_trueOut, cond_br56_trueOut, cond_br47_trueOut, cond_br38_trueOut}),
    .ins_valid ({fork96_outs_1_valid, fork96_outs_0_valid, cond_br308_trueOut_valid, cond_br299_trueOut_valid, cond_br290_trueOut_valid, cond_br281_trueOut_valid, cond_br272_trueOut_valid, cond_br263_trueOut_valid, cond_br254_trueOut_valid, cond_br245_trueOut_valid, cond_br236_trueOut_valid, cond_br227_trueOut_valid, cond_br218_trueOut_valid, cond_br209_trueOut_valid, cond_br200_trueOut_valid, cond_br191_trueOut_valid, cond_br182_trueOut_valid, cond_br173_trueOut_valid, cond_br164_trueOut_valid, cond_br155_trueOut_valid, cond_br146_trueOut_valid, cond_br137_trueOut_valid, cond_br128_trueOut_valid, cond_br119_trueOut_valid, cond_br110_trueOut_valid, cond_br101_trueOut_valid, cond_br92_trueOut_valid, cond_br83_trueOut_valid, cond_br74_trueOut_valid, cond_br65_trueOut_valid, cond_br56_trueOut_valid, cond_br47_trueOut_valid, cond_br38_trueOut_valid}),
    .ins_ready ({fork96_outs_1_ready, fork96_outs_0_ready, cond_br308_trueOut_ready, cond_br299_trueOut_ready, cond_br290_trueOut_ready, cond_br281_trueOut_ready, cond_br272_trueOut_ready, cond_br263_trueOut_ready, cond_br254_trueOut_ready, cond_br245_trueOut_ready, cond_br236_trueOut_ready, cond_br227_trueOut_ready, cond_br218_trueOut_ready, cond_br209_trueOut_ready, cond_br200_trueOut_ready, cond_br191_trueOut_ready, cond_br182_trueOut_ready, cond_br173_trueOut_ready, cond_br164_trueOut_ready, cond_br155_trueOut_ready, cond_br146_trueOut_ready, cond_br137_trueOut_ready, cond_br128_trueOut_ready, cond_br119_trueOut_ready, cond_br110_trueOut_ready, cond_br101_trueOut_ready, cond_br92_trueOut_ready, cond_br83_trueOut_ready, cond_br74_trueOut_ready, cond_br65_trueOut_ready, cond_br56_trueOut_ready, cond_br47_trueOut_ready, cond_br38_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux6_outs),
    .outs_valid (mux6_outs_valid),
    .outs_ready (mux6_outs_ready)
  );

  oehb #(.DATA_TYPE(7)) buffer198(
    .ins (mux6_outs),
    .ins_valid (mux6_outs_valid),
    .ins_ready (mux6_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer198_outs),
    .outs_valid (buffer198_outs_valid),
    .outs_ready (buffer198_outs_ready)
  );

  tehb #(.DATA_TYPE(7)) buffer199(
    .ins (buffer198_outs),
    .ins_valid (buffer198_outs_valid),
    .ins_ready (buffer198_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer199_outs),
    .outs_valid (buffer199_outs_valid),
    .outs_ready (buffer199_outs_ready)
  );

  fork_type #(.SIZE(5), .DATA_TYPE(7)) fork98(
    .ins (buffer199_outs),
    .ins_valid (buffer199_outs_valid),
    .ins_ready (buffer199_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork98_outs_4, fork98_outs_3, fork98_outs_2, fork98_outs_1, fork98_outs_0}),
    .outs_valid ({fork98_outs_4_valid, fork98_outs_3_valid, fork98_outs_2_valid, fork98_outs_1_valid, fork98_outs_0_valid}),
    .outs_ready ({fork98_outs_4_ready, fork98_outs_3_ready, fork98_outs_2_ready, fork98_outs_1_ready, fork98_outs_0_ready})
  );

  control_merge_dataless #(.SIZE(33), .INDEX_TYPE(6)) control_merge31(
    .ins_valid ({fork97_outs_1_valid, fork97_outs_0_valid, cond_br309_trueOut_valid, cond_br300_trueOut_valid, cond_br291_trueOut_valid, cond_br282_trueOut_valid, cond_br273_trueOut_valid, cond_br264_trueOut_valid, cond_br255_trueOut_valid, cond_br246_trueOut_valid, cond_br237_trueOut_valid, cond_br228_trueOut_valid, cond_br219_trueOut_valid, cond_br210_trueOut_valid, cond_br201_trueOut_valid, cond_br192_trueOut_valid, cond_br183_trueOut_valid, cond_br174_trueOut_valid, cond_br165_trueOut_valid, cond_br156_trueOut_valid, cond_br147_trueOut_valid, cond_br138_trueOut_valid, cond_br129_trueOut_valid, cond_br120_trueOut_valid, cond_br111_trueOut_valid, cond_br102_trueOut_valid, cond_br93_trueOut_valid, cond_br84_trueOut_valid, cond_br75_trueOut_valid, cond_br66_trueOut_valid, cond_br57_trueOut_valid, cond_br48_trueOut_valid, cond_br39_trueOut_valid}),
    .ins_ready ({fork97_outs_1_ready, fork97_outs_0_ready, cond_br309_trueOut_ready, cond_br300_trueOut_ready, cond_br291_trueOut_ready, cond_br282_trueOut_ready, cond_br273_trueOut_ready, cond_br264_trueOut_ready, cond_br255_trueOut_ready, cond_br246_trueOut_ready, cond_br237_trueOut_ready, cond_br228_trueOut_ready, cond_br219_trueOut_ready, cond_br210_trueOut_ready, cond_br201_trueOut_ready, cond_br192_trueOut_ready, cond_br183_trueOut_ready, cond_br174_trueOut_ready, cond_br165_trueOut_ready, cond_br156_trueOut_ready, cond_br147_trueOut_ready, cond_br138_trueOut_ready, cond_br129_trueOut_ready, cond_br120_trueOut_ready, cond_br111_trueOut_ready, cond_br102_trueOut_ready, cond_br93_trueOut_ready, cond_br84_trueOut_ready, cond_br75_trueOut_ready, cond_br66_trueOut_ready, cond_br57_trueOut_ready, cond_br48_trueOut_ready, cond_br39_trueOut_ready}),
    .clk (clk),
    .rst (rst),
    .outs_valid (control_merge31_outs_valid),
    .outs_ready (control_merge31_outs_ready),
    .index (control_merge31_index),
    .index_valid (control_merge31_index_valid),
    .index_ready (control_merge31_index_ready)
  );

  fork_type #(.SIZE(7), .DATA_TYPE(6)) fork99(
    .ins (control_merge31_index),
    .ins_valid (control_merge31_index_valid),
    .ins_ready (control_merge31_index_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork99_outs_6, fork99_outs_5, fork99_outs_4, fork99_outs_3, fork99_outs_2, fork99_outs_1, fork99_outs_0}),
    .outs_valid ({fork99_outs_6_valid, fork99_outs_5_valid, fork99_outs_4_valid, fork99_outs_3_valid, fork99_outs_2_valid, fork99_outs_1_valid, fork99_outs_0_valid}),
    .outs_ready ({fork99_outs_6_ready, fork99_outs_5_ready, fork99_outs_4_ready, fork99_outs_3_ready, fork99_outs_2_ready, fork99_outs_1_ready, fork99_outs_0_ready})
  );

  oehb_dataless buffer200(
    .ins_valid (control_merge31_outs_valid),
    .ins_ready (control_merge31_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer200_outs_valid),
    .outs_ready (buffer200_outs_ready)
  );

  tehb_dataless buffer201(
    .ins_valid (buffer200_outs_valid),
    .ins_ready (buffer200_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer201_outs_valid),
    .outs_ready (buffer201_outs_ready)
  );

  sink_dataless sink262(
    .ins_valid (buffer201_outs_valid),
    .ins_ready (buffer201_outs_ready),
    .clk (clk),
    .rst (rst)
  );

  source source33(
    .clk (clk),
    .rst (rst),
    .outs_valid (source33_outs_valid),
    .outs_ready (source33_outs_ready)
  );

  handshake_constant_14 #(.DATA_WIDTH(2)) constant574(
    .ctrl_valid (source33_outs_valid),
    .ctrl_ready (source33_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant574_outs),
    .outs_valid (constant574_outs_valid),
    .outs_ready (constant574_outs_ready)
  );

  fork_type #(.SIZE(5), .DATA_TYPE(2)) fork100(
    .ins (constant574_outs),
    .ins_valid (constant574_outs_valid),
    .ins_ready (constant574_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork100_outs_4, fork100_outs_3, fork100_outs_2, fork100_outs_1, fork100_outs_0}),
    .outs_valid ({fork100_outs_4_valid, fork100_outs_3_valid, fork100_outs_2_valid, fork100_outs_1_valid, fork100_outs_0_valid}),
    .outs_ready ({fork100_outs_4_ready, fork100_outs_3_ready, fork100_outs_2_ready, fork100_outs_1_ready, fork100_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(39)) extsi135(
    .ins (fork100_outs_0),
    .ins_valid (fork100_outs_0_valid),
    .ins_ready (fork100_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi135_outs),
    .outs_valid (extsi135_outs_valid),
    .outs_ready (extsi135_outs_ready)
  );

  extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(35)) extsi136(
    .ins (fork100_outs_1),
    .ins_valid (fork100_outs_1_valid),
    .ins_ready (fork100_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi136_outs),
    .outs_valid (extsi136_outs_valid),
    .outs_ready (extsi136_outs_ready)
  );

  extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(29)) extsi137(
    .ins (fork100_outs_2),
    .ins_valid (fork100_outs_2_valid),
    .ins_ready (fork100_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi137_outs),
    .outs_valid (extsi137_outs_valid),
    .outs_ready (extsi137_outs_ready)
  );

  extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(24)) extsi138(
    .ins (fork100_outs_3),
    .ins_valid (fork100_outs_3_valid),
    .ins_ready (fork100_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi138_outs),
    .outs_valid (extsi138_outs_valid),
    .outs_ready (extsi138_outs_ready)
  );

  extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(19)) extsi139(
    .ins (fork100_outs_4),
    .ins_valid (fork100_outs_4_valid),
    .ins_ready (fork100_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi139_outs),
    .outs_valid (extsi139_outs_valid),
    .outs_ready (extsi139_outs_ready)
  );

  source source38(
    .clk (clk),
    .rst (rst),
    .outs_valid (source38_outs_valid),
    .outs_ready (source38_outs_ready)
  );

  handshake_constant_35 #(.DATA_WIDTH(4)) constant575(
    .ctrl_valid (source38_outs_valid),
    .ctrl_ready (source38_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant575_outs),
    .outs_valid (constant575_outs_valid),
    .outs_ready (constant575_outs_ready)
  );

  extui #(.INPUT_TYPE(4), .OUTPUT_TYPE(12)) extui0(
    .ins (constant575_outs),
    .ins_valid (constant575_outs_valid),
    .ins_ready (constant575_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extui0_outs),
    .outs_valid (extui0_outs_valid),
    .outs_ready (extui0_outs_ready)
  );

  trunci #(.INPUT_TYPE(7), .OUTPUT_TYPE(6)) trunci1(
    .ins (fork98_outs_4),
    .ins_valid (fork98_outs_4_valid),
    .ins_ready (fork98_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci1_outs),
    .outs_valid (trunci1_outs_valid),
    .outs_ready (trunci1_outs_ready)
  );

  oehb #(.DATA_TYPE(12)) buffer196(
    .ins (mux5_outs),
    .ins_valid (mux5_outs_valid),
    .ins_ready (mux5_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer196_outs),
    .outs_valid (buffer196_outs_valid),
    .outs_ready (buffer196_outs_ready)
  );

  tehb #(.DATA_TYPE(12)) buffer197(
    .ins (buffer196_outs),
    .ins_valid (buffer196_outs_valid),
    .ins_ready (buffer196_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer197_outs),
    .outs_valid (buffer197_outs_valid),
    .outs_ready (buffer197_outs_ready)
  );

  extsi #(.INPUT_TYPE(12), .OUTPUT_TYPE(18)) extsi0(
    .ins (buffer197_outs),
    .ins_valid (buffer197_outs_valid),
    .ins_ready (buffer197_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi0_outs),
    .outs_valid (extsi0_outs_valid),
    .outs_ready (extsi0_outs_ready)
  );

  extsi #(.INPUT_TYPE(6), .OUTPUT_TYPE(18)) extsi1(
    .ins (trunci1_outs),
    .ins_valid (trunci1_outs_valid),
    .ins_ready (trunci1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi1_outs),
    .outs_valid (extsi1_outs_valid),
    .outs_ready (extsi1_outs_ready)
  );

  muli #(.DATA_TYPE(18)) muli0(
    .lhs (extsi0_outs),
    .lhs_valid (extsi0_outs_valid),
    .lhs_ready (extsi0_outs_ready),
    .rhs (extsi1_outs),
    .rhs_valid (extsi1_outs_valid),
    .rhs_ready (extsi1_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli0_result),
    .result_valid (muli0_result_valid),
    .result_ready (muli0_result_ready)
  );

  oehb #(.DATA_TYPE(17)) buffer194(
    .ins (mux4_outs),
    .ins_valid (mux4_outs_valid),
    .ins_ready (mux4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer194_outs),
    .outs_valid (buffer194_outs_valid),
    .outs_ready (buffer194_outs_ready)
  );

  tehb #(.DATA_TYPE(17)) buffer195(
    .ins (buffer194_outs),
    .ins_valid (buffer194_outs_valid),
    .ins_ready (buffer194_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer195_outs),
    .outs_valid (buffer195_outs_valid),
    .outs_ready (buffer195_outs_ready)
  );

  extsi #(.INPUT_TYPE(17), .OUTPUT_TYPE(19)) extsi3(
    .ins (buffer195_outs),
    .ins_valid (buffer195_outs_valid),
    .ins_ready (buffer195_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi3_outs),
    .outs_valid (extsi3_outs_valid),
    .outs_ready (extsi3_outs_ready)
  );

  shli #(.DATA_TYPE(19)) shli0(
    .lhs (extsi3_outs),
    .lhs_valid (extsi3_outs_valid),
    .lhs_ready (extsi3_outs_ready),
    .rhs (extsi139_outs),
    .rhs_valid (extsi139_outs_valid),
    .rhs_ready (extsi139_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli0_result),
    .result_valid (shli0_result_valid),
    .result_ready (shli0_result_ready)
  );

  trunci #(.INPUT_TYPE(19), .OUTPUT_TYPE(18)) trunci14(
    .ins (shli0_result),
    .ins_valid (shli0_result_valid),
    .ins_ready (shli0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci14_outs),
    .outs_valid (trunci14_outs_valid),
    .outs_ready (trunci14_outs_ready)
  );

  addi #(.DATA_TYPE(18)) addi0(
    .lhs (muli0_result),
    .lhs_valid (muli0_result_valid),
    .lhs_ready (muli0_result_ready),
    .rhs (trunci14_outs),
    .rhs_valid (trunci14_outs_valid),
    .rhs_ready (trunci14_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi0_result),
    .result_valid (addi0_result_valid),
    .result_ready (addi0_result_ready)
  );

  extsi #(.INPUT_TYPE(18), .OUTPUT_TYPE(25)) extsi4(
    .ins (addi0_result),
    .ins_valid (addi0_result_valid),
    .ins_ready (addi0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi4_outs),
    .outs_valid (extsi4_outs_valid),
    .outs_ready (extsi4_outs_ready)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(25)) extsi5(
    .ins (fork98_outs_0),
    .ins_valid (fork98_outs_0_valid),
    .ins_ready (fork98_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi5_outs),
    .outs_valid (extsi5_outs_valid),
    .outs_ready (extsi5_outs_ready)
  );

  muli #(.DATA_TYPE(25)) muli1(
    .lhs (extsi4_outs),
    .lhs_valid (extsi4_outs_valid),
    .lhs_ready (extsi4_outs_ready),
    .rhs (extsi5_outs),
    .rhs_valid (extsi5_outs_valid),
    .rhs_ready (extsi5_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli1_result),
    .result_valid (muli1_result_valid),
    .result_ready (muli1_result_ready)
  );

  trunci #(.INPUT_TYPE(25), .OUTPUT_TYPE(23)) trunci4(
    .ins (muli1_result),
    .ins_valid (muli1_result_valid),
    .ins_ready (muli1_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci4_outs),
    .outs_valid (trunci4_outs_valid),
    .outs_ready (trunci4_outs_ready)
  );

  oehb #(.DATA_TYPE(22)) buffer192(
    .ins (mux3_outs),
    .ins_valid (mux3_outs_valid),
    .ins_ready (mux3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer192_outs),
    .outs_valid (buffer192_outs_valid),
    .outs_ready (buffer192_outs_ready)
  );

  tehb #(.DATA_TYPE(22)) buffer193(
    .ins (buffer192_outs),
    .ins_valid (buffer192_outs_valid),
    .ins_ready (buffer192_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer193_outs),
    .outs_valid (buffer193_outs_valid),
    .outs_ready (buffer193_outs_ready)
  );

  extsi #(.INPUT_TYPE(22), .OUTPUT_TYPE(24)) extsi7(
    .ins (buffer193_outs),
    .ins_valid (buffer193_outs_valid),
    .ins_ready (buffer193_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi7_outs),
    .outs_valid (extsi7_outs_valid),
    .outs_ready (extsi7_outs_ready)
  );

  shli #(.DATA_TYPE(24)) shli1(
    .lhs (extsi7_outs),
    .lhs_valid (extsi7_outs_valid),
    .lhs_ready (extsi7_outs_ready),
    .rhs (extsi138_outs),
    .rhs_valid (extsi138_outs_valid),
    .rhs_ready (extsi138_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli1_result),
    .result_valid (shli1_result_valid),
    .result_ready (shli1_result_ready)
  );

  trunci #(.INPUT_TYPE(24), .OUTPUT_TYPE(23)) trunci15(
    .ins (shli1_result),
    .ins_valid (shli1_result_valid),
    .ins_ready (shli1_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci15_outs),
    .outs_valid (trunci15_outs_valid),
    .outs_ready (trunci15_outs_ready)
  );

  addi #(.DATA_TYPE(23)) addi1(
    .lhs (trunci4_outs),
    .lhs_valid (trunci4_outs_valid),
    .lhs_ready (trunci4_outs_ready),
    .rhs (trunci15_outs),
    .rhs_valid (trunci15_outs_valid),
    .rhs_ready (trunci15_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi1_result),
    .result_valid (addi1_result_valid),
    .result_ready (addi1_result_ready)
  );

  extsi #(.INPUT_TYPE(23), .OUTPUT_TYPE(30)) extsi8(
    .ins (addi1_result),
    .ins_valid (addi1_result_valid),
    .ins_ready (addi1_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi8_outs),
    .outs_valid (extsi8_outs_valid),
    .outs_ready (extsi8_outs_ready)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(30)) extsi9(
    .ins (fork98_outs_1),
    .ins_valid (fork98_outs_1_valid),
    .ins_ready (fork98_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi9_outs),
    .outs_valid (extsi9_outs_valid),
    .outs_ready (extsi9_outs_ready)
  );

  muli #(.DATA_TYPE(30)) muli2(
    .lhs (extsi8_outs),
    .lhs_valid (extsi8_outs_valid),
    .lhs_ready (extsi8_outs_ready),
    .rhs (extsi9_outs),
    .rhs_valid (extsi9_outs_valid),
    .rhs_ready (extsi9_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli2_result),
    .result_valid (muli2_result_valid),
    .result_ready (muli2_result_ready)
  );

  trunci #(.INPUT_TYPE(30), .OUTPUT_TYPE(28)) trunci6(
    .ins (muli2_result),
    .ins_valid (muli2_result_valid),
    .ins_ready (muli2_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci6_outs),
    .outs_valid (trunci6_outs_valid),
    .outs_ready (trunci6_outs_ready)
  );

  oehb #(.DATA_TYPE(27)) buffer190(
    .ins (mux2_outs),
    .ins_valid (mux2_outs_valid),
    .ins_ready (mux2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer190_outs),
    .outs_valid (buffer190_outs_valid),
    .outs_ready (buffer190_outs_ready)
  );

  tehb #(.DATA_TYPE(27)) buffer191(
    .ins (buffer190_outs),
    .ins_valid (buffer190_outs_valid),
    .ins_ready (buffer190_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer191_outs),
    .outs_valid (buffer191_outs_valid),
    .outs_ready (buffer191_outs_ready)
  );

  extsi #(.INPUT_TYPE(27), .OUTPUT_TYPE(29)) extsi11(
    .ins (buffer191_outs),
    .ins_valid (buffer191_outs_valid),
    .ins_ready (buffer191_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi11_outs),
    .outs_valid (extsi11_outs_valid),
    .outs_ready (extsi11_outs_ready)
  );

  shli #(.DATA_TYPE(29)) shli2(
    .lhs (extsi11_outs),
    .lhs_valid (extsi11_outs_valid),
    .lhs_ready (extsi11_outs_ready),
    .rhs (extsi137_outs),
    .rhs_valid (extsi137_outs_valid),
    .rhs_ready (extsi137_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli2_result),
    .result_valid (shli2_result_valid),
    .result_ready (shli2_result_ready)
  );

  trunci #(.INPUT_TYPE(29), .OUTPUT_TYPE(28)) trunci16(
    .ins (shli2_result),
    .ins_valid (shli2_result_valid),
    .ins_ready (shli2_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci16_outs),
    .outs_valid (trunci16_outs_valid),
    .outs_ready (trunci16_outs_ready)
  );

  addi #(.DATA_TYPE(28)) addi2(
    .lhs (trunci6_outs),
    .lhs_valid (trunci6_outs_valid),
    .lhs_ready (trunci6_outs_ready),
    .rhs (trunci16_outs),
    .rhs_valid (trunci16_outs_valid),
    .rhs_ready (trunci16_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi2_result),
    .result_valid (addi2_result_valid),
    .result_ready (addi2_result_ready)
  );

  extsi #(.INPUT_TYPE(28), .OUTPUT_TYPE(35)) extsi12(
    .ins (addi2_result),
    .ins_valid (addi2_result_valid),
    .ins_ready (addi2_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi12_outs),
    .outs_valid (extsi12_outs_valid),
    .outs_ready (extsi12_outs_ready)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(35)) extsi13(
    .ins (fork98_outs_2),
    .ins_valid (fork98_outs_2_valid),
    .ins_ready (fork98_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi13_outs),
    .outs_valid (extsi13_outs_valid),
    .outs_ready (extsi13_outs_ready)
  );

  muli #(.DATA_TYPE(35)) muli3(
    .lhs (extsi12_outs),
    .lhs_valid (extsi12_outs_valid),
    .lhs_ready (extsi12_outs_ready),
    .rhs (extsi13_outs),
    .rhs_valid (extsi13_outs_valid),
    .rhs_ready (extsi13_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli3_result),
    .result_valid (muli3_result_valid),
    .result_ready (muli3_result_ready)
  );

  trunci #(.INPUT_TYPE(35), .OUTPUT_TYPE(34)) trunci8(
    .ins (muli3_result),
    .ins_valid (muli3_result_valid),
    .ins_ready (muli3_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci8_outs),
    .outs_valid (trunci8_outs_valid),
    .outs_ready (trunci8_outs_ready)
  );

  oehb #(.DATA_TYPE(33)) buffer188(
    .ins (mux1_outs),
    .ins_valid (mux1_outs_valid),
    .ins_ready (mux1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer188_outs),
    .outs_valid (buffer188_outs_valid),
    .outs_ready (buffer188_outs_ready)
  );

  tehb #(.DATA_TYPE(33)) buffer189(
    .ins (buffer188_outs),
    .ins_valid (buffer188_outs_valid),
    .ins_ready (buffer188_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer189_outs),
    .outs_valid (buffer189_outs_valid),
    .outs_ready (buffer189_outs_ready)
  );

  extsi #(.INPUT_TYPE(33), .OUTPUT_TYPE(35)) extsi15(
    .ins (buffer189_outs),
    .ins_valid (buffer189_outs_valid),
    .ins_ready (buffer189_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi15_outs),
    .outs_valid (extsi15_outs_valid),
    .outs_ready (extsi15_outs_ready)
  );

  shli #(.DATA_TYPE(35)) shli3(
    .lhs (extsi15_outs),
    .lhs_valid (extsi15_outs_valid),
    .lhs_ready (extsi15_outs_ready),
    .rhs (extsi136_outs),
    .rhs_valid (extsi136_outs_valid),
    .rhs_ready (extsi136_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli3_result),
    .result_valid (shli3_result_valid),
    .result_ready (shli3_result_ready)
  );

  trunci #(.INPUT_TYPE(35), .OUTPUT_TYPE(34)) trunci17(
    .ins (shli3_result),
    .ins_valid (shli3_result_valid),
    .ins_ready (shli3_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci17_outs),
    .outs_valid (trunci17_outs_valid),
    .outs_ready (trunci17_outs_ready)
  );

  addi #(.DATA_TYPE(34)) addi3(
    .lhs (trunci8_outs),
    .lhs_valid (trunci8_outs_valid),
    .lhs_ready (trunci8_outs_ready),
    .rhs (trunci17_outs),
    .rhs_valid (trunci17_outs_valid),
    .rhs_ready (trunci17_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi3_result),
    .result_valid (addi3_result_valid),
    .result_ready (addi3_result_ready)
  );

  extsi #(.INPUT_TYPE(34), .OUTPUT_TYPE(41)) extsi16(
    .ins (addi3_result),
    .ins_valid (addi3_result_valid),
    .ins_ready (addi3_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi16_outs),
    .outs_valid (extsi16_outs_valid),
    .outs_ready (extsi16_outs_ready)
  );

  extsi #(.INPUT_TYPE(7), .OUTPUT_TYPE(41)) extsi17(
    .ins (fork98_outs_3),
    .ins_valid (fork98_outs_3_valid),
    .ins_ready (fork98_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi17_outs),
    .outs_valid (extsi17_outs_valid),
    .outs_ready (extsi17_outs_ready)
  );

  muli #(.DATA_TYPE(41)) muli4(
    .lhs (extsi16_outs),
    .lhs_valid (extsi16_outs_valid),
    .lhs_ready (extsi16_outs_ready),
    .rhs (extsi17_outs),
    .rhs_valid (extsi17_outs_valid),
    .rhs_ready (extsi17_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli4_result),
    .result_valid (muli4_result_valid),
    .result_ready (muli4_result_ready)
  );

  trunci #(.INPUT_TYPE(41), .OUTPUT_TYPE(12)) trunci18(
    .ins (muli4_result),
    .ins_valid (muli4_result_valid),
    .ins_ready (muli4_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci18_outs),
    .outs_valid (trunci18_outs_valid),
    .outs_ready (trunci18_outs_ready)
  );

  oehb #(.DATA_TYPE(37)) buffer186(
    .ins (mux0_outs),
    .ins_valid (mux0_outs_valid),
    .ins_ready (mux0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer186_outs),
    .outs_valid (buffer186_outs_valid),
    .outs_ready (buffer186_outs_ready)
  );

  tehb #(.DATA_TYPE(37)) buffer187(
    .ins (buffer186_outs),
    .ins_valid (buffer186_outs_valid),
    .ins_ready (buffer186_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer187_outs),
    .outs_valid (buffer187_outs_valid),
    .outs_ready (buffer187_outs_ready)
  );

  extsi #(.INPUT_TYPE(37), .OUTPUT_TYPE(39)) extsi19(
    .ins (buffer187_outs),
    .ins_valid (buffer187_outs_valid),
    .ins_ready (buffer187_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi19_outs),
    .outs_valid (extsi19_outs_valid),
    .outs_ready (extsi19_outs_ready)
  );

  shli #(.DATA_TYPE(39)) shli4(
    .lhs (extsi19_outs),
    .lhs_valid (extsi19_outs_valid),
    .lhs_ready (extsi19_outs_ready),
    .rhs (extsi135_outs),
    .rhs_valid (extsi135_outs_valid),
    .rhs_ready (extsi135_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shli4_result),
    .result_valid (shli4_result_valid),
    .result_ready (shli4_result_ready)
  );

  trunci #(.INPUT_TYPE(39), .OUTPUT_TYPE(12)) trunci19(
    .ins (shli4_result),
    .ins_valid (shli4_result_valid),
    .ins_ready (shli4_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci19_outs),
    .outs_valid (trunci19_outs_valid),
    .outs_ready (trunci19_outs_ready)
  );

  addi #(.DATA_TYPE(12)) addi4(
    .lhs (trunci18_outs),
    .lhs_valid (trunci18_outs_valid),
    .lhs_ready (trunci18_outs_ready),
    .rhs (trunci19_outs),
    .rhs_valid (trunci19_outs_valid),
    .rhs_ready (trunci19_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi4_result),
    .result_valid (addi4_result_valid),
    .result_ready (addi4_result_ready)
  );

  shrsi #(.DATA_TYPE(12)) shrsi0(
    .lhs (addi4_result),
    .lhs_valid (addi4_result_valid),
    .lhs_ready (addi4_result_ready),
    .rhs (extui0_outs),
    .rhs_valid (extui0_outs_valid),
    .rhs_ready (extui0_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shrsi0_result),
    .result_valid (shrsi0_result_valid),
    .result_ready (shrsi0_result_ready)
  );

  trunci #(.INPUT_TYPE(12), .OUTPUT_TYPE(8)) trunci12(
    .ins (shrsi0_result),
    .ins_valid (shrsi0_result_valid),
    .ins_ready (shrsi0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci12_outs),
    .outs_valid (trunci12_outs_valid),
    .outs_ready (trunci12_outs_ready)
  );

endmodule
